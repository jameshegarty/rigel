module incif_1uint32(input CLK, input CE, input [32:0] process_input, output [31:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [31:0] unnamedcast12465USEDMULTIPLEcast = (process_input[31:0]);
  assign process_output = (((process_input[32]))?({(unnamedcast12465USEDMULTIPLEcast+(32'd1))}):(unnamedcast12465USEDMULTIPLEcast));
  // function: process pure=true delay=0
endmodule

module RegBy_incif_1uint32_CEtrue_initnil(input CLK, input set_valid, input CE, input [31:0] set_inp, input setby_valid, input setby_inp, output [31:0] SETBY_OUTPUT, output [31:0] GET_OUTPUT);
parameter INSTANCE_NAME="INST";
  reg [31:0] R;
  wire [31:0] regby_inner_process_output;
  always @(posedge CLK) begin if(set_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(setby_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,set_valid})+({4'b0,setby_valid})) > 5'd1) begin $display("error, function 'set' on instance 'R' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [32:0] unnamedcallArbitrate12497USEDMULTIPLEcallArbitrate = {(set_valid||setby_valid),((set_valid)?(set_inp):(regby_inner_process_output))};
    always @ (posedge CLK) begin if ((unnamedcallArbitrate12497USEDMULTIPLEcallArbitrate[32]) && CE) begin R <= (unnamedcallArbitrate12497USEDMULTIPLEcallArbitrate[31:0]); end end
  assign SETBY_OUTPUT = regby_inner_process_output;
  assign GET_OUTPUT = R;
  // function: set pure=false ONLY WIRE
  // function: setby pure=false ONLY WIRE
  // function: get pure=true ONLY WIRE
  incif_1uint32 #(.INSTANCE_NAME("regby_inner")) regby_inner(.CLK(CLK), .CE(CE), .process_input({setby_inp,R}), .process_output(regby_inner_process_output));
endmodule

module Underflow_Auint8_8_1__count38400_cycles154624_toosoonnil_UStrue(input CLK, input ready_downstream, output ready, input reset, input [64:0] process_input, output [64:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire [31:0] cycleCount_GET_OUTPUT;
  wire unnamedbinop13129USEDMULTIPLEbinop = {((cycleCount_GET_OUTPUT)>((32'd154624)))};
  assign ready = {(ready_downstream||unnamedbinop13129USEDMULTIPLEbinop)};
  wire unnamedbinop13131USEDMULTIPLEbinop = {({(ready_downstream||reset)}||unnamedbinop13129USEDMULTIPLEbinop)};
  wire [31:0] outputCount_GET_OUTPUT;
  wire unnamedcast13123USEDMULTIPLEcast = (process_input[64]);
  wire unnamedunary13151USEDMULTIPLEunary = {(~reset)};
  wire [31:0] outputCount_SETBY_OUTPUT;
  wire [31:0] cycleCount_SETBY_OUTPUT;
  assign process_output = {{({({(unnamedbinop13129USEDMULTIPLEbinop&&{((outputCount_GET_OUTPUT)<((32'd38400)))})}||{({(~unnamedbinop13129USEDMULTIPLEbinop)}&&unnamedcast13123USEDMULTIPLEcast)})}&&unnamedunary13151USEDMULTIPLEunary)},((unnamedbinop13129USEDMULTIPLEbinop)?((64'd3735928559)):((process_input[63:0])))};
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  RegBy_incif_1uint32_CEtrue_initnil #(.INSTANCE_NAME("outputCount")) outputCount(.CLK(CLK), .set_valid(reset), .CE(unnamedbinop13131USEDMULTIPLEbinop), .set_inp((32'd0)), .setby_valid(unnamedunary13151USEDMULTIPLEunary), .setby_inp({(ready_downstream&&{(unnamedcast13123USEDMULTIPLEcast||unnamedbinop13129USEDMULTIPLEbinop)})}), .SETBY_OUTPUT(outputCount_SETBY_OUTPUT), .GET_OUTPUT(outputCount_GET_OUTPUT));
  RegBy_incif_1uint32_CEtrue_initnil #(.INSTANCE_NAME("cycleCount")) cycleCount(.CLK(CLK), .set_valid(reset), .CE((1'd1)), .set_inp((32'd0)), .setby_valid(unnamedunary13151USEDMULTIPLEunary), .setby_inp((1'd1)), .SETBY_OUTPUT(cycleCount_SETBY_OUTPUT), .GET_OUTPUT(cycleCount_GET_OUTPUT));
endmodule

module incif_wrap127_incnil(input CLK, input CE, input [8:0] process_input, output [7:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [7:0] unnamedcast384USEDMULTIPLEcast = (process_input[7:0]);
  assign process_output = (((process_input[8]))?((({(unnamedcast384USEDMULTIPLEcast==(8'd127))})?((8'd0)):({(unnamedcast384USEDMULTIPLEcast+(8'd1))}))):(unnamedcast384USEDMULTIPLEcast));
  // function: process pure=true delay=0
endmodule

module RegBy_incif_wrap127_incnil_CEtrue_initnil(input CLK, input set_valid, input CE, input [7:0] set_inp, input setby_valid, input setby_inp, output [7:0] SETBY_OUTPUT, output [7:0] GET_OUTPUT);
parameter INSTANCE_NAME="INST";
  reg [7:0] R;
  wire [7:0] regby_inner_process_output;
  always @(posedge CLK) begin if(set_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(setby_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,set_valid})+({4'b0,setby_valid})) > 5'd1) begin $display("error, function 'set' on instance 'R' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [8:0] unnamedcallArbitrate435USEDMULTIPLEcallArbitrate = {(set_valid||setby_valid),((set_valid)?(set_inp):(regby_inner_process_output))};
    always @ (posedge CLK) begin if ((unnamedcallArbitrate435USEDMULTIPLEcallArbitrate[8]) && CE) begin R <= (unnamedcallArbitrate435USEDMULTIPLEcallArbitrate[7:0]); end end
  assign SETBY_OUTPUT = regby_inner_process_output;
  assign GET_OUTPUT = R;
  // function: set pure=false ONLY WIRE
  // function: setby pure=false ONLY WIRE
  // function: get pure=true ONLY WIRE
  incif_wrap127_incnil #(.INSTANCE_NAME("regby_inner")) regby_inner(.CLK(CLK), .CE(CE), .process_input({setby_inp,R}), .process_output(regby_inner_process_output));
endmodule

module fifo_uint8_8_1_(input CLK, input popFront_valid, input CE_pop, output [63:0] popFront, output [7:0] size, input pushBackReset_valid, input CE_push, output ready, input pushBack_valid, input [63:0] pushBack_input, input popFrontReset_valid, output hasData);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(popFront_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'popFront'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(pushBackReset_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'pushBackReset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(pushBack_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'pushBack'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(popFrontReset_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'popFrontReset'", INSTANCE_NAME);  end end
  wire [7:0] readAddr_GET_OUTPUT;
  wire [6:0] unnamedcast791USEDMULTIPLEcast = readAddr_GET_OUTPUT[6:0];
  wire fifo1_READ_OUTPUT;
  wire fifo2_READ_OUTPUT;
  wire fifo3_READ_OUTPUT;
  wire fifo4_READ_OUTPUT;
  wire fifo5_READ_OUTPUT;
  wire fifo6_READ_OUTPUT;
  wire fifo7_READ_OUTPUT;
  wire fifo8_READ_OUTPUT;
  wire fifo9_READ_OUTPUT;
  wire fifo10_READ_OUTPUT;
  wire fifo11_READ_OUTPUT;
  wire fifo12_READ_OUTPUT;
  wire fifo13_READ_OUTPUT;
  wire fifo14_READ_OUTPUT;
  wire fifo15_READ_OUTPUT;
  wire fifo16_READ_OUTPUT;
  wire fifo17_READ_OUTPUT;
  wire fifo18_READ_OUTPUT;
  wire fifo19_READ_OUTPUT;
  wire fifo20_READ_OUTPUT;
  wire fifo21_READ_OUTPUT;
  wire fifo22_READ_OUTPUT;
  wire fifo23_READ_OUTPUT;
  wire fifo24_READ_OUTPUT;
  wire fifo25_READ_OUTPUT;
  wire fifo26_READ_OUTPUT;
  wire fifo27_READ_OUTPUT;
  wire fifo28_READ_OUTPUT;
  wire fifo29_READ_OUTPUT;
  wire fifo30_READ_OUTPUT;
  wire fifo31_READ_OUTPUT;
  wire fifo32_READ_OUTPUT;
  wire fifo33_READ_OUTPUT;
  wire fifo34_READ_OUTPUT;
  wire fifo35_READ_OUTPUT;
  wire fifo36_READ_OUTPUT;
  wire fifo37_READ_OUTPUT;
  wire fifo38_READ_OUTPUT;
  wire fifo39_READ_OUTPUT;
  wire fifo40_READ_OUTPUT;
  wire fifo41_READ_OUTPUT;
  wire fifo42_READ_OUTPUT;
  wire fifo43_READ_OUTPUT;
  wire fifo44_READ_OUTPUT;
  wire fifo45_READ_OUTPUT;
  wire fifo46_READ_OUTPUT;
  wire fifo47_READ_OUTPUT;
  wire fifo48_READ_OUTPUT;
  wire fifo49_READ_OUTPUT;
  wire fifo50_READ_OUTPUT;
  wire fifo51_READ_OUTPUT;
  wire fifo52_READ_OUTPUT;
  wire fifo53_READ_OUTPUT;
  wire fifo54_READ_OUTPUT;
  wire fifo55_READ_OUTPUT;
  wire fifo56_READ_OUTPUT;
  wire fifo57_READ_OUTPUT;
  wire fifo58_READ_OUTPUT;
  wire fifo59_READ_OUTPUT;
  wire fifo60_READ_OUTPUT;
  wire fifo61_READ_OUTPUT;
  wire fifo62_READ_OUTPUT;
  wire fifo63_READ_OUTPUT;
  wire fifo64_READ_OUTPUT;
  wire [7:0] writeAddr_GET_OUTPUT;
  wire unnamedunary458USEDMULTIPLEunary = {(~{(writeAddr_GET_OUTPUT==readAddr_GET_OUTPUT)})};
  always @(posedge CLK) begin if(unnamedunary458USEDMULTIPLEunary == 1'b0 && popFront_valid==1'b1 && CE_pop==1'b1) begin $display("%s: attempting to pop from an empty fifo",INSTANCE_NAME);$finish();  end end
  wire [7:0] readAddr_SETBY_OUTPUT;
  assign popFront = {fifo64_READ_OUTPUT,fifo63_READ_OUTPUT,fifo62_READ_OUTPUT,fifo61_READ_OUTPUT,fifo60_READ_OUTPUT,fifo59_READ_OUTPUT,fifo58_READ_OUTPUT,fifo57_READ_OUTPUT,fifo56_READ_OUTPUT,fifo55_READ_OUTPUT,fifo54_READ_OUTPUT,fifo53_READ_OUTPUT,fifo52_READ_OUTPUT,fifo51_READ_OUTPUT,fifo50_READ_OUTPUT,fifo49_READ_OUTPUT,fifo48_READ_OUTPUT,fifo47_READ_OUTPUT,fifo46_READ_OUTPUT,fifo45_READ_OUTPUT,fifo44_READ_OUTPUT,fifo43_READ_OUTPUT,fifo42_READ_OUTPUT,fifo41_READ_OUTPUT,fifo40_READ_OUTPUT,fifo39_READ_OUTPUT,fifo38_READ_OUTPUT,fifo37_READ_OUTPUT,fifo36_READ_OUTPUT,fifo35_READ_OUTPUT,fifo34_READ_OUTPUT,fifo33_READ_OUTPUT,fifo32_READ_OUTPUT,fifo31_READ_OUTPUT,fifo30_READ_OUTPUT,fifo29_READ_OUTPUT,fifo28_READ_OUTPUT,fifo27_READ_OUTPUT,fifo26_READ_OUTPUT,fifo25_READ_OUTPUT,fifo24_READ_OUTPUT,fifo23_READ_OUTPUT,fifo22_READ_OUTPUT,fifo21_READ_OUTPUT,fifo20_READ_OUTPUT,fifo19_READ_OUTPUT,fifo18_READ_OUTPUT,fifo17_READ_OUTPUT,fifo16_READ_OUTPUT,fifo15_READ_OUTPUT,fifo14_READ_OUTPUT,fifo13_READ_OUTPUT,fifo12_READ_OUTPUT,fifo11_READ_OUTPUT,fifo10_READ_OUTPUT,fifo9_READ_OUTPUT,fifo8_READ_OUTPUT,fifo7_READ_OUTPUT,fifo6_READ_OUTPUT,fifo5_READ_OUTPUT,fifo4_READ_OUTPUT,fifo3_READ_OUTPUT,fifo2_READ_OUTPUT,fifo1_READ_OUTPUT};
  wire [7:0] unnamedselect449USEDMULTIPLEselect = (({((writeAddr_GET_OUTPUT)<(readAddr_GET_OUTPUT))})?({({((8'd128)-readAddr_GET_OUTPUT)}+writeAddr_GET_OUTPUT)}):({(writeAddr_GET_OUTPUT-readAddr_GET_OUTPUT)}));
  assign size = unnamedselect449USEDMULTIPLEselect;
  reg readyReg;
    always @ (posedge CLK) begin readyReg <= {((unnamedselect449USEDMULTIPLEselect)<((8'd125)))}; end
  assign ready = readyReg;
  always @(posedge CLK) begin if({((unnamedselect449USEDMULTIPLEselect)<((8'd126)))} == 1'b0 && pushBack_valid==1'b1 && CE_push==1'b1) begin $display("%s: attempting to push to a full fifo",INSTANCE_NAME);$finish();  end end
  wire [7:0] writeAddr_SETBY_OUTPUT;
  wire [6:0] unnamedcast466USEDMULTIPLEcast = writeAddr_GET_OUTPUT[6:0];
  assign hasData = unnamedunary458USEDMULTIPLEunary;
  // function: popFront pure=false delay=0
  // function: size pure=true delay=0
  // function: pushBackReset pure=false delay=0
  // function: ready pure=true delay=0
  // function: pushBack pure=false delay=0
  // function: popFrontReset pure=false delay=0
  // function: hasData pure=true delay=0
  RegBy_incif_wrap127_incnil_CEtrue_initnil #(.INSTANCE_NAME("writeAddr")) writeAddr(.CLK(CLK), .set_valid(pushBackReset_valid), .CE(CE_push), .set_inp((8'd0)), .setby_valid(pushBack_valid), .setby_inp((1'd1)), .SETBY_OUTPUT(writeAddr_SETBY_OUTPUT), .GET_OUTPUT(writeAddr_GET_OUTPUT));
  RegBy_incif_wrap127_incnil_CEtrue_initnil #(.INSTANCE_NAME("readAddr")) readAddr(.CLK(CLK), .set_valid(popFrontReset_valid), .CE(CE_pop), .set_inp((8'd0)), .setby_valid(popFront_valid), .setby_inp((1'd1)), .SETBY_OUTPUT(readAddr_SETBY_OUTPUT), .GET_OUTPUT(readAddr_GET_OUTPUT));
  wire [7:0] fifo1_writeInput = {pushBack_input[0:0],unnamedcast466USEDMULTIPLEcast};
wire fifo1_writeOut;
RAM128X1D fifo1  (
  .WCLK(CLK),
  .D(fifo1_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo1_writeOut),
  .DPO(fifo1_READ_OUTPUT),
  .A(fifo1_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo2_writeInput = {pushBack_input[1:1],unnamedcast466USEDMULTIPLEcast};
wire fifo2_writeOut;
RAM128X1D fifo2  (
  .WCLK(CLK),
  .D(fifo2_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo2_writeOut),
  .DPO(fifo2_READ_OUTPUT),
  .A(fifo2_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo3_writeInput = {pushBack_input[2:2],unnamedcast466USEDMULTIPLEcast};
wire fifo3_writeOut;
RAM128X1D fifo3  (
  .WCLK(CLK),
  .D(fifo3_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo3_writeOut),
  .DPO(fifo3_READ_OUTPUT),
  .A(fifo3_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo4_writeInput = {pushBack_input[3:3],unnamedcast466USEDMULTIPLEcast};
wire fifo4_writeOut;
RAM128X1D fifo4  (
  .WCLK(CLK),
  .D(fifo4_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo4_writeOut),
  .DPO(fifo4_READ_OUTPUT),
  .A(fifo4_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo5_writeInput = {pushBack_input[4:4],unnamedcast466USEDMULTIPLEcast};
wire fifo5_writeOut;
RAM128X1D fifo5  (
  .WCLK(CLK),
  .D(fifo5_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo5_writeOut),
  .DPO(fifo5_READ_OUTPUT),
  .A(fifo5_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo6_writeInput = {pushBack_input[5:5],unnamedcast466USEDMULTIPLEcast};
wire fifo6_writeOut;
RAM128X1D fifo6  (
  .WCLK(CLK),
  .D(fifo6_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo6_writeOut),
  .DPO(fifo6_READ_OUTPUT),
  .A(fifo6_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo7_writeInput = {pushBack_input[6:6],unnamedcast466USEDMULTIPLEcast};
wire fifo7_writeOut;
RAM128X1D fifo7  (
  .WCLK(CLK),
  .D(fifo7_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo7_writeOut),
  .DPO(fifo7_READ_OUTPUT),
  .A(fifo7_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo8_writeInput = {pushBack_input[7:7],unnamedcast466USEDMULTIPLEcast};
wire fifo8_writeOut;
RAM128X1D fifo8  (
  .WCLK(CLK),
  .D(fifo8_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo8_writeOut),
  .DPO(fifo8_READ_OUTPUT),
  .A(fifo8_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo9_writeInput = {pushBack_input[8:8],unnamedcast466USEDMULTIPLEcast};
wire fifo9_writeOut;
RAM128X1D fifo9  (
  .WCLK(CLK),
  .D(fifo9_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo9_writeOut),
  .DPO(fifo9_READ_OUTPUT),
  .A(fifo9_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo10_writeInput = {pushBack_input[9:9],unnamedcast466USEDMULTIPLEcast};
wire fifo10_writeOut;
RAM128X1D fifo10  (
  .WCLK(CLK),
  .D(fifo10_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo10_writeOut),
  .DPO(fifo10_READ_OUTPUT),
  .A(fifo10_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo11_writeInput = {pushBack_input[10:10],unnamedcast466USEDMULTIPLEcast};
wire fifo11_writeOut;
RAM128X1D fifo11  (
  .WCLK(CLK),
  .D(fifo11_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo11_writeOut),
  .DPO(fifo11_READ_OUTPUT),
  .A(fifo11_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo12_writeInput = {pushBack_input[11:11],unnamedcast466USEDMULTIPLEcast};
wire fifo12_writeOut;
RAM128X1D fifo12  (
  .WCLK(CLK),
  .D(fifo12_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo12_writeOut),
  .DPO(fifo12_READ_OUTPUT),
  .A(fifo12_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo13_writeInput = {pushBack_input[12:12],unnamedcast466USEDMULTIPLEcast};
wire fifo13_writeOut;
RAM128X1D fifo13  (
  .WCLK(CLK),
  .D(fifo13_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo13_writeOut),
  .DPO(fifo13_READ_OUTPUT),
  .A(fifo13_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo14_writeInput = {pushBack_input[13:13],unnamedcast466USEDMULTIPLEcast};
wire fifo14_writeOut;
RAM128X1D fifo14  (
  .WCLK(CLK),
  .D(fifo14_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo14_writeOut),
  .DPO(fifo14_READ_OUTPUT),
  .A(fifo14_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo15_writeInput = {pushBack_input[14:14],unnamedcast466USEDMULTIPLEcast};
wire fifo15_writeOut;
RAM128X1D fifo15  (
  .WCLK(CLK),
  .D(fifo15_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo15_writeOut),
  .DPO(fifo15_READ_OUTPUT),
  .A(fifo15_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo16_writeInput = {pushBack_input[15:15],unnamedcast466USEDMULTIPLEcast};
wire fifo16_writeOut;
RAM128X1D fifo16  (
  .WCLK(CLK),
  .D(fifo16_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo16_writeOut),
  .DPO(fifo16_READ_OUTPUT),
  .A(fifo16_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo17_writeInput = {pushBack_input[16:16],unnamedcast466USEDMULTIPLEcast};
wire fifo17_writeOut;
RAM128X1D fifo17  (
  .WCLK(CLK),
  .D(fifo17_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo17_writeOut),
  .DPO(fifo17_READ_OUTPUT),
  .A(fifo17_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo18_writeInput = {pushBack_input[17:17],unnamedcast466USEDMULTIPLEcast};
wire fifo18_writeOut;
RAM128X1D fifo18  (
  .WCLK(CLK),
  .D(fifo18_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo18_writeOut),
  .DPO(fifo18_READ_OUTPUT),
  .A(fifo18_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo19_writeInput = {pushBack_input[18:18],unnamedcast466USEDMULTIPLEcast};
wire fifo19_writeOut;
RAM128X1D fifo19  (
  .WCLK(CLK),
  .D(fifo19_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo19_writeOut),
  .DPO(fifo19_READ_OUTPUT),
  .A(fifo19_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo20_writeInput = {pushBack_input[19:19],unnamedcast466USEDMULTIPLEcast};
wire fifo20_writeOut;
RAM128X1D fifo20  (
  .WCLK(CLK),
  .D(fifo20_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo20_writeOut),
  .DPO(fifo20_READ_OUTPUT),
  .A(fifo20_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo21_writeInput = {pushBack_input[20:20],unnamedcast466USEDMULTIPLEcast};
wire fifo21_writeOut;
RAM128X1D fifo21  (
  .WCLK(CLK),
  .D(fifo21_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo21_writeOut),
  .DPO(fifo21_READ_OUTPUT),
  .A(fifo21_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo22_writeInput = {pushBack_input[21:21],unnamedcast466USEDMULTIPLEcast};
wire fifo22_writeOut;
RAM128X1D fifo22  (
  .WCLK(CLK),
  .D(fifo22_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo22_writeOut),
  .DPO(fifo22_READ_OUTPUT),
  .A(fifo22_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo23_writeInput = {pushBack_input[22:22],unnamedcast466USEDMULTIPLEcast};
wire fifo23_writeOut;
RAM128X1D fifo23  (
  .WCLK(CLK),
  .D(fifo23_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo23_writeOut),
  .DPO(fifo23_READ_OUTPUT),
  .A(fifo23_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo24_writeInput = {pushBack_input[23:23],unnamedcast466USEDMULTIPLEcast};
wire fifo24_writeOut;
RAM128X1D fifo24  (
  .WCLK(CLK),
  .D(fifo24_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo24_writeOut),
  .DPO(fifo24_READ_OUTPUT),
  .A(fifo24_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo25_writeInput = {pushBack_input[24:24],unnamedcast466USEDMULTIPLEcast};
wire fifo25_writeOut;
RAM128X1D fifo25  (
  .WCLK(CLK),
  .D(fifo25_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo25_writeOut),
  .DPO(fifo25_READ_OUTPUT),
  .A(fifo25_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo26_writeInput = {pushBack_input[25:25],unnamedcast466USEDMULTIPLEcast};
wire fifo26_writeOut;
RAM128X1D fifo26  (
  .WCLK(CLK),
  .D(fifo26_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo26_writeOut),
  .DPO(fifo26_READ_OUTPUT),
  .A(fifo26_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo27_writeInput = {pushBack_input[26:26],unnamedcast466USEDMULTIPLEcast};
wire fifo27_writeOut;
RAM128X1D fifo27  (
  .WCLK(CLK),
  .D(fifo27_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo27_writeOut),
  .DPO(fifo27_READ_OUTPUT),
  .A(fifo27_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo28_writeInput = {pushBack_input[27:27],unnamedcast466USEDMULTIPLEcast};
wire fifo28_writeOut;
RAM128X1D fifo28  (
  .WCLK(CLK),
  .D(fifo28_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo28_writeOut),
  .DPO(fifo28_READ_OUTPUT),
  .A(fifo28_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo29_writeInput = {pushBack_input[28:28],unnamedcast466USEDMULTIPLEcast};
wire fifo29_writeOut;
RAM128X1D fifo29  (
  .WCLK(CLK),
  .D(fifo29_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo29_writeOut),
  .DPO(fifo29_READ_OUTPUT),
  .A(fifo29_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo30_writeInput = {pushBack_input[29:29],unnamedcast466USEDMULTIPLEcast};
wire fifo30_writeOut;
RAM128X1D fifo30  (
  .WCLK(CLK),
  .D(fifo30_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo30_writeOut),
  .DPO(fifo30_READ_OUTPUT),
  .A(fifo30_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo31_writeInput = {pushBack_input[30:30],unnamedcast466USEDMULTIPLEcast};
wire fifo31_writeOut;
RAM128X1D fifo31  (
  .WCLK(CLK),
  .D(fifo31_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo31_writeOut),
  .DPO(fifo31_READ_OUTPUT),
  .A(fifo31_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo32_writeInput = {pushBack_input[31:31],unnamedcast466USEDMULTIPLEcast};
wire fifo32_writeOut;
RAM128X1D fifo32  (
  .WCLK(CLK),
  .D(fifo32_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo32_writeOut),
  .DPO(fifo32_READ_OUTPUT),
  .A(fifo32_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo33_writeInput = {pushBack_input[32:32],unnamedcast466USEDMULTIPLEcast};
wire fifo33_writeOut;
RAM128X1D fifo33  (
  .WCLK(CLK),
  .D(fifo33_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo33_writeOut),
  .DPO(fifo33_READ_OUTPUT),
  .A(fifo33_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo34_writeInput = {pushBack_input[33:33],unnamedcast466USEDMULTIPLEcast};
wire fifo34_writeOut;
RAM128X1D fifo34  (
  .WCLK(CLK),
  .D(fifo34_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo34_writeOut),
  .DPO(fifo34_READ_OUTPUT),
  .A(fifo34_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo35_writeInput = {pushBack_input[34:34],unnamedcast466USEDMULTIPLEcast};
wire fifo35_writeOut;
RAM128X1D fifo35  (
  .WCLK(CLK),
  .D(fifo35_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo35_writeOut),
  .DPO(fifo35_READ_OUTPUT),
  .A(fifo35_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo36_writeInput = {pushBack_input[35:35],unnamedcast466USEDMULTIPLEcast};
wire fifo36_writeOut;
RAM128X1D fifo36  (
  .WCLK(CLK),
  .D(fifo36_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo36_writeOut),
  .DPO(fifo36_READ_OUTPUT),
  .A(fifo36_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo37_writeInput = {pushBack_input[36:36],unnamedcast466USEDMULTIPLEcast};
wire fifo37_writeOut;
RAM128X1D fifo37  (
  .WCLK(CLK),
  .D(fifo37_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo37_writeOut),
  .DPO(fifo37_READ_OUTPUT),
  .A(fifo37_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo38_writeInput = {pushBack_input[37:37],unnamedcast466USEDMULTIPLEcast};
wire fifo38_writeOut;
RAM128X1D fifo38  (
  .WCLK(CLK),
  .D(fifo38_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo38_writeOut),
  .DPO(fifo38_READ_OUTPUT),
  .A(fifo38_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo39_writeInput = {pushBack_input[38:38],unnamedcast466USEDMULTIPLEcast};
wire fifo39_writeOut;
RAM128X1D fifo39  (
  .WCLK(CLK),
  .D(fifo39_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo39_writeOut),
  .DPO(fifo39_READ_OUTPUT),
  .A(fifo39_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo40_writeInput = {pushBack_input[39:39],unnamedcast466USEDMULTIPLEcast};
wire fifo40_writeOut;
RAM128X1D fifo40  (
  .WCLK(CLK),
  .D(fifo40_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo40_writeOut),
  .DPO(fifo40_READ_OUTPUT),
  .A(fifo40_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo41_writeInput = {pushBack_input[40:40],unnamedcast466USEDMULTIPLEcast};
wire fifo41_writeOut;
RAM128X1D fifo41  (
  .WCLK(CLK),
  .D(fifo41_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo41_writeOut),
  .DPO(fifo41_READ_OUTPUT),
  .A(fifo41_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo42_writeInput = {pushBack_input[41:41],unnamedcast466USEDMULTIPLEcast};
wire fifo42_writeOut;
RAM128X1D fifo42  (
  .WCLK(CLK),
  .D(fifo42_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo42_writeOut),
  .DPO(fifo42_READ_OUTPUT),
  .A(fifo42_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo43_writeInput = {pushBack_input[42:42],unnamedcast466USEDMULTIPLEcast};
wire fifo43_writeOut;
RAM128X1D fifo43  (
  .WCLK(CLK),
  .D(fifo43_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo43_writeOut),
  .DPO(fifo43_READ_OUTPUT),
  .A(fifo43_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo44_writeInput = {pushBack_input[43:43],unnamedcast466USEDMULTIPLEcast};
wire fifo44_writeOut;
RAM128X1D fifo44  (
  .WCLK(CLK),
  .D(fifo44_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo44_writeOut),
  .DPO(fifo44_READ_OUTPUT),
  .A(fifo44_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo45_writeInput = {pushBack_input[44:44],unnamedcast466USEDMULTIPLEcast};
wire fifo45_writeOut;
RAM128X1D fifo45  (
  .WCLK(CLK),
  .D(fifo45_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo45_writeOut),
  .DPO(fifo45_READ_OUTPUT),
  .A(fifo45_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo46_writeInput = {pushBack_input[45:45],unnamedcast466USEDMULTIPLEcast};
wire fifo46_writeOut;
RAM128X1D fifo46  (
  .WCLK(CLK),
  .D(fifo46_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo46_writeOut),
  .DPO(fifo46_READ_OUTPUT),
  .A(fifo46_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo47_writeInput = {pushBack_input[46:46],unnamedcast466USEDMULTIPLEcast};
wire fifo47_writeOut;
RAM128X1D fifo47  (
  .WCLK(CLK),
  .D(fifo47_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo47_writeOut),
  .DPO(fifo47_READ_OUTPUT),
  .A(fifo47_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo48_writeInput = {pushBack_input[47:47],unnamedcast466USEDMULTIPLEcast};
wire fifo48_writeOut;
RAM128X1D fifo48  (
  .WCLK(CLK),
  .D(fifo48_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo48_writeOut),
  .DPO(fifo48_READ_OUTPUT),
  .A(fifo48_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo49_writeInput = {pushBack_input[48:48],unnamedcast466USEDMULTIPLEcast};
wire fifo49_writeOut;
RAM128X1D fifo49  (
  .WCLK(CLK),
  .D(fifo49_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo49_writeOut),
  .DPO(fifo49_READ_OUTPUT),
  .A(fifo49_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo50_writeInput = {pushBack_input[49:49],unnamedcast466USEDMULTIPLEcast};
wire fifo50_writeOut;
RAM128X1D fifo50  (
  .WCLK(CLK),
  .D(fifo50_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo50_writeOut),
  .DPO(fifo50_READ_OUTPUT),
  .A(fifo50_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo51_writeInput = {pushBack_input[50:50],unnamedcast466USEDMULTIPLEcast};
wire fifo51_writeOut;
RAM128X1D fifo51  (
  .WCLK(CLK),
  .D(fifo51_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo51_writeOut),
  .DPO(fifo51_READ_OUTPUT),
  .A(fifo51_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo52_writeInput = {pushBack_input[51:51],unnamedcast466USEDMULTIPLEcast};
wire fifo52_writeOut;
RAM128X1D fifo52  (
  .WCLK(CLK),
  .D(fifo52_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo52_writeOut),
  .DPO(fifo52_READ_OUTPUT),
  .A(fifo52_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo53_writeInput = {pushBack_input[52:52],unnamedcast466USEDMULTIPLEcast};
wire fifo53_writeOut;
RAM128X1D fifo53  (
  .WCLK(CLK),
  .D(fifo53_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo53_writeOut),
  .DPO(fifo53_READ_OUTPUT),
  .A(fifo53_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo54_writeInput = {pushBack_input[53:53],unnamedcast466USEDMULTIPLEcast};
wire fifo54_writeOut;
RAM128X1D fifo54  (
  .WCLK(CLK),
  .D(fifo54_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo54_writeOut),
  .DPO(fifo54_READ_OUTPUT),
  .A(fifo54_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo55_writeInput = {pushBack_input[54:54],unnamedcast466USEDMULTIPLEcast};
wire fifo55_writeOut;
RAM128X1D fifo55  (
  .WCLK(CLK),
  .D(fifo55_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo55_writeOut),
  .DPO(fifo55_READ_OUTPUT),
  .A(fifo55_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo56_writeInput = {pushBack_input[55:55],unnamedcast466USEDMULTIPLEcast};
wire fifo56_writeOut;
RAM128X1D fifo56  (
  .WCLK(CLK),
  .D(fifo56_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo56_writeOut),
  .DPO(fifo56_READ_OUTPUT),
  .A(fifo56_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo57_writeInput = {pushBack_input[56:56],unnamedcast466USEDMULTIPLEcast};
wire fifo57_writeOut;
RAM128X1D fifo57  (
  .WCLK(CLK),
  .D(fifo57_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo57_writeOut),
  .DPO(fifo57_READ_OUTPUT),
  .A(fifo57_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo58_writeInput = {pushBack_input[57:57],unnamedcast466USEDMULTIPLEcast};
wire fifo58_writeOut;
RAM128X1D fifo58  (
  .WCLK(CLK),
  .D(fifo58_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo58_writeOut),
  .DPO(fifo58_READ_OUTPUT),
  .A(fifo58_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo59_writeInput = {pushBack_input[58:58],unnamedcast466USEDMULTIPLEcast};
wire fifo59_writeOut;
RAM128X1D fifo59  (
  .WCLK(CLK),
  .D(fifo59_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo59_writeOut),
  .DPO(fifo59_READ_OUTPUT),
  .A(fifo59_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo60_writeInput = {pushBack_input[59:59],unnamedcast466USEDMULTIPLEcast};
wire fifo60_writeOut;
RAM128X1D fifo60  (
  .WCLK(CLK),
  .D(fifo60_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo60_writeOut),
  .DPO(fifo60_READ_OUTPUT),
  .A(fifo60_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo61_writeInput = {pushBack_input[60:60],unnamedcast466USEDMULTIPLEcast};
wire fifo61_writeOut;
RAM128X1D fifo61  (
  .WCLK(CLK),
  .D(fifo61_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo61_writeOut),
  .DPO(fifo61_READ_OUTPUT),
  .A(fifo61_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo62_writeInput = {pushBack_input[61:61],unnamedcast466USEDMULTIPLEcast};
wire fifo62_writeOut;
RAM128X1D fifo62  (
  .WCLK(CLK),
  .D(fifo62_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo62_writeOut),
  .DPO(fifo62_READ_OUTPUT),
  .A(fifo62_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo63_writeInput = {pushBack_input[62:62],unnamedcast466USEDMULTIPLEcast};
wire fifo63_writeOut;
RAM128X1D fifo63  (
  .WCLK(CLK),
  .D(fifo63_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo63_writeOut),
  .DPO(fifo63_READ_OUTPUT),
  .A(fifo63_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

  wire [7:0] fifo64_writeInput = {pushBack_input[63:63],unnamedcast466USEDMULTIPLEcast};
wire fifo64_writeOut;
RAM128X1D fifo64  (
  .WCLK(CLK),
  .D(fifo64_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo64_writeOut),
  .DPO(fifo64_READ_OUTPUT),
  .A(fifo64_writeInput[6:0]),
  .DPRA(unnamedcast791USEDMULTIPLEcast));

endmodule

module fifo_128_uint8_8_1_(input CLK, input load_valid, input load_CE, output [64:0] load_output, input store_reset_valid, input store_CE, output store_ready, input load_reset_valid, input store_valid, input [63:0] store_input);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(load_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_reset_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(load_reset_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store'", INSTANCE_NAME);  end end
  wire FIFO_hasData;
  wire [63:0] FIFO_popFront;
  assign load_output = {FIFO_hasData,FIFO_popFront};
  wire FIFO_ready;
  assign store_ready = FIFO_ready;
  // function: load pure=false delay=0
  // function: store_reset pure=false delay=0
  // function: store_ready pure=true delay=0
  // function: load_reset pure=false delay=0
  // function: store pure=false delay=0
  fifo_uint8_8_1_ #(.INSTANCE_NAME("FIFO")) FIFO(.CLK(CLK), .popFront_valid({(FIFO_hasData&&load_valid)}), .CE_pop(load_CE), .popFront(FIFO_popFront), .size(FIFO_size), .pushBackReset_valid(store_reset_valid), .CE_push(store_CE), .ready(FIFO_ready), .pushBack_valid(store_valid), .pushBack_input(store_input), .popFrontReset_valid(load_reset_valid), .hasData(FIFO_hasData));
endmodule

module LiftDecimate_fifo_128_uint8_8_1_(input CLK, input load_valid, input load_CE, input load_input, output [64:0] load_output, input store_reset_valid, input store_CE, output store_ready, output load_ready, input load_reset, input store_valid, input [63:0] store_input);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(load_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_reset_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(load_reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store'", INSTANCE_NAME);  end end
  wire unnamedcast1890USEDMULTIPLEcast = load_input;
  wire [64:0] LiftDecimate_inner_fifo_128_uint8_8_1__load_output;
  reg [63:0] unnamedcast1893_delay1_validunnamednull0_CEload_CE;  always @ (posedge CLK) begin if (load_CE) begin unnamedcast1893_delay1_validunnamednull0_CEload_CE <= (LiftDecimate_inner_fifo_128_uint8_8_1__load_output[63:0]); end end
  reg unnamedbinop1898_delay1_validunnamednull0_CEload_CE;  always @ (posedge CLK) begin if (load_CE) begin unnamedbinop1898_delay1_validunnamednull0_CEload_CE <= {((LiftDecimate_inner_fifo_128_uint8_8_1__load_output[64])&&unnamedcast1890USEDMULTIPLEcast)}; end end
  assign load_output = {unnamedbinop1898_delay1_validunnamednull0_CEload_CE,unnamedcast1893_delay1_validunnamednull0_CEload_CE};
  wire LiftDecimate_inner_fifo_128_uint8_8_1__store_ready;
  assign store_ready = LiftDecimate_inner_fifo_128_uint8_8_1__store_ready;
  assign load_ready = (1'd1);
  // function: load pure=false delay=1
  // function: store_reset pure=false delay=0
  // function: store_ready pure=true delay=0
  // function: load_ready pure=true delay=0
  // function: load_reset pure=false delay=0
  // function: store pure=false delay=0
  fifo_128_uint8_8_1_ #(.INSTANCE_NAME("LiftDecimate_inner_fifo_128_uint8_8_1_")) LiftDecimate_inner_fifo_128_uint8_8_1_(.CLK(CLK), .load_valid({(unnamedcast1890USEDMULTIPLEcast&&load_valid)}), .load_CE(load_CE), .load_output(LiftDecimate_inner_fifo_128_uint8_8_1__load_output), .store_reset_valid(store_reset_valid), .store_CE(store_CE), .store_ready(LiftDecimate_inner_fifo_128_uint8_8_1__store_ready), .load_reset_valid(load_reset), .store_valid(store_valid), .store_input(store_input));
endmodule

module RunIffReady_LiftDecimate_fifo_128_uint8_8_1_(input CLK, input load_valid, input load_CE, input load_input, output [64:0] load_output, input store_reset, input CE, output store_ready, output load_ready, input load_reset, input store_valid, input [64:0] store_input, output store_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(load_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(load_reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store'", INSTANCE_NAME);  end end
  wire [64:0] RunIffReady_inner_load_output;
  assign load_output = RunIffReady_inner_load_output;
  wire RunIffReady_inner_store_ready;
  assign store_ready = RunIffReady_inner_store_ready;
  wire RunIffReady_inner_load_ready;
  assign load_ready = RunIffReady_inner_load_ready;
  wire unnamedbinop1969USEDMULTIPLEbinop = {({(RunIffReady_inner_store_ready&&(store_input[64]))}&&store_valid)};
  assign store_output = {unnamedbinop1969USEDMULTIPLEbinop};
  // function: load pure=false delay=1
  // function: store_reset pure=false delay=0
  // function: store_ready pure=true delay=0
  // function: load_ready pure=true delay=0
  // function: load_reset pure=false delay=0
  // function: store pure=false delay=0
  LiftDecimate_fifo_128_uint8_8_1_ #(.INSTANCE_NAME("RunIffReady_inner")) RunIffReady_inner(.CLK(CLK), .load_valid(load_valid), .load_CE(load_CE), .load_input(load_input), .load_output(RunIffReady_inner_load_output), .store_reset_valid(store_reset), .store_CE(CE), .store_ready(RunIffReady_inner_store_ready), .load_ready(RunIffReady_inner_load_ready), .load_reset(load_reset), .store_valid(unnamedbinop1969USEDMULTIPLEbinop), .store_input((store_input[63:0])));
endmodule

module ShiftRegister_1_CEtrue_TY1(input CLK, input pushPop_valid, input CE, input sr_input, output pushPop_out, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'pushPop'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  reg SR1;
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR1' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR1' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR1' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate352USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(sr_input):((1'd0)))};
    always @ (posedge CLK) begin if ((unnamedcallArbitrate352USEDMULTIPLEcallArbitrate[1]) && CE) begin SR1 <= (unnamedcallArbitrate352USEDMULTIPLEcallArbitrate[0]); end end
  assign pushPop_out = SR1;
  // function: pushPop pure=false delay=0
  // function: reset pure=false delay=0
endmodule

module ShiftRegister_0_CEtrue_TY1(input CLK, input CE, input sr_input, output pushPop_out);
parameter INSTANCE_NAME="INST";
  assign pushPop_out = sr_input;
  // function: pushPop pure=true delay=0
  // function: reset pure=true delay=0
endmodule

module LiftHandshake_RunIffReady_LiftDecimate_fifo_128_uint8_8_1_(input CLK, input load_input, output [64:0] load_output, input store_reset, input store_ready_downstream, output store_ready, input load_ready_downstream, output load_ready, input load_reset, input [64:0] store_input, output store_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire unnamedunary2006USEDMULTIPLEunary = {(~load_reset)};
  wire unnamedbinop2005USEDMULTIPLEbinop = {(load_reset||load_ready_downstream)};
  wire [64:0] inner_RunIffReady_LiftDecimate_fifo_128_uint8_8_1__load_output;
  wire load_validBitDelay_RunIffReady_LiftDecimate_fifo_128_uint8_8_1__pushPop_out;
  wire [64:0] unnamedtuple2016USEDMULTIPLEtuple = {{((inner_RunIffReady_LiftDecimate_fifo_128_uint8_8_1__load_output[64])&&load_validBitDelay_RunIffReady_LiftDecimate_fifo_128_uint8_8_1__pushPop_out)},(inner_RunIffReady_LiftDecimate_fifo_128_uint8_8_1__load_output[63:0])};
  always @(posedge CLK) begin if({(~{((unnamedtuple2016USEDMULTIPLEtuple[64])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: output valid bit should not be X!",INSTANCE_NAME); end end
  always @(posedge CLK) begin if({(~{(load_input===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign load_output = unnamedtuple2016USEDMULTIPLEtuple;
  wire unnamedbinop2034USEDMULTIPLEbinop = {(store_reset||store_ready_downstream)};
  wire inner_RunIffReady_LiftDecimate_fifo_128_uint8_8_1__store_ready;
  assign store_ready = {(inner_RunIffReady_LiftDecimate_fifo_128_uint8_8_1__store_ready&&store_ready_downstream)};
  wire inner_RunIffReady_LiftDecimate_fifo_128_uint8_8_1__load_ready;
  assign load_ready = {(inner_RunIffReady_LiftDecimate_fifo_128_uint8_8_1__load_ready&&load_ready_downstream)};
  wire unnamedunary2035USEDMULTIPLEunary = {(~store_reset)};
  wire [0:0] inner_RunIffReady_LiftDecimate_fifo_128_uint8_8_1__store_output;
  wire store_validBitDelay_RunIffReady_LiftDecimate_fifo_128_uint8_8_1__pushPop_out;
  wire [0:0] unnamedtuple2049USEDMULTIPLEtuple = {{(inner_RunIffReady_LiftDecimate_fifo_128_uint8_8_1__store_output&&store_validBitDelay_RunIffReady_LiftDecimate_fifo_128_uint8_8_1__pushPop_out)}};
  always @(posedge CLK) begin if({(~{(unnamedtuple2049USEDMULTIPLEtuple===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: output valid bit should not be X!",INSTANCE_NAME); end end
  always @(posedge CLK) begin if({(~{((store_input[64])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign store_output = unnamedtuple2049USEDMULTIPLEtuple;
  // function: load pure=false ONLY WIRE
  // function: store_reset pure=false ONLY WIRE
  // function: store_ready pure=true ONLY WIRE
  // function: load_ready pure=true ONLY WIRE
  // function: load_reset pure=false ONLY WIRE
  // function: store pure=false ONLY WIRE
  RunIffReady_LiftDecimate_fifo_128_uint8_8_1_ #(.INSTANCE_NAME("inner_RunIffReady_LiftDecimate_fifo_128_uint8_8_1_")) inner_RunIffReady_LiftDecimate_fifo_128_uint8_8_1_(.CLK(CLK), .load_valid(unnamedunary2006USEDMULTIPLEunary), .load_CE(unnamedbinop2005USEDMULTIPLEbinop), .load_input(load_input), .load_output(inner_RunIffReady_LiftDecimate_fifo_128_uint8_8_1__load_output), .store_reset(store_reset), .CE(unnamedbinop2034USEDMULTIPLEbinop), .store_ready(inner_RunIffReady_LiftDecimate_fifo_128_uint8_8_1__store_ready), .load_ready(inner_RunIffReady_LiftDecimate_fifo_128_uint8_8_1__load_ready), .load_reset(load_reset), .store_valid(unnamedunary2035USEDMULTIPLEunary), .store_input(store_input), .store_output(inner_RunIffReady_LiftDecimate_fifo_128_uint8_8_1__store_output));
  ShiftRegister_1_CEtrue_TY1 #(.INSTANCE_NAME("load_validBitDelay_RunIffReady_LiftDecimate_fifo_128_uint8_8_1_")) load_validBitDelay_RunIffReady_LiftDecimate_fifo_128_uint8_8_1_(.CLK(CLK), .pushPop_valid(unnamedunary2006USEDMULTIPLEunary), .CE(unnamedbinop2005USEDMULTIPLEbinop), .sr_input((1'd1)), .pushPop_out(load_validBitDelay_RunIffReady_LiftDecimate_fifo_128_uint8_8_1__pushPop_out), .reset(load_reset));
  ShiftRegister_0_CEtrue_TY1 #(.INSTANCE_NAME("store_validBitDelay_RunIffReady_LiftDecimate_fifo_128_uint8_8_1_")) store_validBitDelay_RunIffReady_LiftDecimate_fifo_128_uint8_8_1_(.CLK(CLK), .CE(unnamedbinop2034USEDMULTIPLEbinop), .sr_input((1'd1)), .pushPop_out(store_validBitDelay_RunIffReady_LiftDecimate_fifo_128_uint8_8_1__pushPop_out));
endmodule

module fifo_uint8_4_1__8_1_(input CLK, input popFront_valid, input CE_pop, output [255:0] popFront, output [7:0] size, input pushBackReset_valid, input CE_push, output ready, input pushBack_valid, input [255:0] pushBack_input, input popFrontReset_valid, output hasData);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(popFront_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'popFront'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(pushBackReset_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'pushBackReset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(pushBack_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'pushBack'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(popFrontReset_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'popFrontReset'", INSTANCE_NAME);  end end
  wire [7:0] readAddr_GET_OUTPUT;
  wire [6:0] unnamedcast7992USEDMULTIPLEcast = readAddr_GET_OUTPUT[6:0];
  wire fifo1_READ_OUTPUT;
  wire fifo2_READ_OUTPUT;
  wire fifo3_READ_OUTPUT;
  wire fifo4_READ_OUTPUT;
  wire fifo5_READ_OUTPUT;
  wire fifo6_READ_OUTPUT;
  wire fifo7_READ_OUTPUT;
  wire fifo8_READ_OUTPUT;
  wire fifo9_READ_OUTPUT;
  wire fifo10_READ_OUTPUT;
  wire fifo11_READ_OUTPUT;
  wire fifo12_READ_OUTPUT;
  wire fifo13_READ_OUTPUT;
  wire fifo14_READ_OUTPUT;
  wire fifo15_READ_OUTPUT;
  wire fifo16_READ_OUTPUT;
  wire fifo17_READ_OUTPUT;
  wire fifo18_READ_OUTPUT;
  wire fifo19_READ_OUTPUT;
  wire fifo20_READ_OUTPUT;
  wire fifo21_READ_OUTPUT;
  wire fifo22_READ_OUTPUT;
  wire fifo23_READ_OUTPUT;
  wire fifo24_READ_OUTPUT;
  wire fifo25_READ_OUTPUT;
  wire fifo26_READ_OUTPUT;
  wire fifo27_READ_OUTPUT;
  wire fifo28_READ_OUTPUT;
  wire fifo29_READ_OUTPUT;
  wire fifo30_READ_OUTPUT;
  wire fifo31_READ_OUTPUT;
  wire fifo32_READ_OUTPUT;
  wire fifo33_READ_OUTPUT;
  wire fifo34_READ_OUTPUT;
  wire fifo35_READ_OUTPUT;
  wire fifo36_READ_OUTPUT;
  wire fifo37_READ_OUTPUT;
  wire fifo38_READ_OUTPUT;
  wire fifo39_READ_OUTPUT;
  wire fifo40_READ_OUTPUT;
  wire fifo41_READ_OUTPUT;
  wire fifo42_READ_OUTPUT;
  wire fifo43_READ_OUTPUT;
  wire fifo44_READ_OUTPUT;
  wire fifo45_READ_OUTPUT;
  wire fifo46_READ_OUTPUT;
  wire fifo47_READ_OUTPUT;
  wire fifo48_READ_OUTPUT;
  wire fifo49_READ_OUTPUT;
  wire fifo50_READ_OUTPUT;
  wire fifo51_READ_OUTPUT;
  wire fifo52_READ_OUTPUT;
  wire fifo53_READ_OUTPUT;
  wire fifo54_READ_OUTPUT;
  wire fifo55_READ_OUTPUT;
  wire fifo56_READ_OUTPUT;
  wire fifo57_READ_OUTPUT;
  wire fifo58_READ_OUTPUT;
  wire fifo59_READ_OUTPUT;
  wire fifo60_READ_OUTPUT;
  wire fifo61_READ_OUTPUT;
  wire fifo62_READ_OUTPUT;
  wire fifo63_READ_OUTPUT;
  wire fifo64_READ_OUTPUT;
  wire fifo65_READ_OUTPUT;
  wire fifo66_READ_OUTPUT;
  wire fifo67_READ_OUTPUT;
  wire fifo68_READ_OUTPUT;
  wire fifo69_READ_OUTPUT;
  wire fifo70_READ_OUTPUT;
  wire fifo71_READ_OUTPUT;
  wire fifo72_READ_OUTPUT;
  wire fifo73_READ_OUTPUT;
  wire fifo74_READ_OUTPUT;
  wire fifo75_READ_OUTPUT;
  wire fifo76_READ_OUTPUT;
  wire fifo77_READ_OUTPUT;
  wire fifo78_READ_OUTPUT;
  wire fifo79_READ_OUTPUT;
  wire fifo80_READ_OUTPUT;
  wire fifo81_READ_OUTPUT;
  wire fifo82_READ_OUTPUT;
  wire fifo83_READ_OUTPUT;
  wire fifo84_READ_OUTPUT;
  wire fifo85_READ_OUTPUT;
  wire fifo86_READ_OUTPUT;
  wire fifo87_READ_OUTPUT;
  wire fifo88_READ_OUTPUT;
  wire fifo89_READ_OUTPUT;
  wire fifo90_READ_OUTPUT;
  wire fifo91_READ_OUTPUT;
  wire fifo92_READ_OUTPUT;
  wire fifo93_READ_OUTPUT;
  wire fifo94_READ_OUTPUT;
  wire fifo95_READ_OUTPUT;
  wire fifo96_READ_OUTPUT;
  wire fifo97_READ_OUTPUT;
  wire fifo98_READ_OUTPUT;
  wire fifo99_READ_OUTPUT;
  wire fifo100_READ_OUTPUT;
  wire fifo101_READ_OUTPUT;
  wire fifo102_READ_OUTPUT;
  wire fifo103_READ_OUTPUT;
  wire fifo104_READ_OUTPUT;
  wire fifo105_READ_OUTPUT;
  wire fifo106_READ_OUTPUT;
  wire fifo107_READ_OUTPUT;
  wire fifo108_READ_OUTPUT;
  wire fifo109_READ_OUTPUT;
  wire fifo110_READ_OUTPUT;
  wire fifo111_READ_OUTPUT;
  wire fifo112_READ_OUTPUT;
  wire fifo113_READ_OUTPUT;
  wire fifo114_READ_OUTPUT;
  wire fifo115_READ_OUTPUT;
  wire fifo116_READ_OUTPUT;
  wire fifo117_READ_OUTPUT;
  wire fifo118_READ_OUTPUT;
  wire fifo119_READ_OUTPUT;
  wire fifo120_READ_OUTPUT;
  wire fifo121_READ_OUTPUT;
  wire fifo122_READ_OUTPUT;
  wire fifo123_READ_OUTPUT;
  wire fifo124_READ_OUTPUT;
  wire fifo125_READ_OUTPUT;
  wire fifo126_READ_OUTPUT;
  wire fifo127_READ_OUTPUT;
  wire fifo128_READ_OUTPUT;
  wire fifo129_READ_OUTPUT;
  wire fifo130_READ_OUTPUT;
  wire fifo131_READ_OUTPUT;
  wire fifo132_READ_OUTPUT;
  wire fifo133_READ_OUTPUT;
  wire fifo134_READ_OUTPUT;
  wire fifo135_READ_OUTPUT;
  wire fifo136_READ_OUTPUT;
  wire fifo137_READ_OUTPUT;
  wire fifo138_READ_OUTPUT;
  wire fifo139_READ_OUTPUT;
  wire fifo140_READ_OUTPUT;
  wire fifo141_READ_OUTPUT;
  wire fifo142_READ_OUTPUT;
  wire fifo143_READ_OUTPUT;
  wire fifo144_READ_OUTPUT;
  wire fifo145_READ_OUTPUT;
  wire fifo146_READ_OUTPUT;
  wire fifo147_READ_OUTPUT;
  wire fifo148_READ_OUTPUT;
  wire fifo149_READ_OUTPUT;
  wire fifo150_READ_OUTPUT;
  wire fifo151_READ_OUTPUT;
  wire fifo152_READ_OUTPUT;
  wire fifo153_READ_OUTPUT;
  wire fifo154_READ_OUTPUT;
  wire fifo155_READ_OUTPUT;
  wire fifo156_READ_OUTPUT;
  wire fifo157_READ_OUTPUT;
  wire fifo158_READ_OUTPUT;
  wire fifo159_READ_OUTPUT;
  wire fifo160_READ_OUTPUT;
  wire fifo161_READ_OUTPUT;
  wire fifo162_READ_OUTPUT;
  wire fifo163_READ_OUTPUT;
  wire fifo164_READ_OUTPUT;
  wire fifo165_READ_OUTPUT;
  wire fifo166_READ_OUTPUT;
  wire fifo167_READ_OUTPUT;
  wire fifo168_READ_OUTPUT;
  wire fifo169_READ_OUTPUT;
  wire fifo170_READ_OUTPUT;
  wire fifo171_READ_OUTPUT;
  wire fifo172_READ_OUTPUT;
  wire fifo173_READ_OUTPUT;
  wire fifo174_READ_OUTPUT;
  wire fifo175_READ_OUTPUT;
  wire fifo176_READ_OUTPUT;
  wire fifo177_READ_OUTPUT;
  wire fifo178_READ_OUTPUT;
  wire fifo179_READ_OUTPUT;
  wire fifo180_READ_OUTPUT;
  wire fifo181_READ_OUTPUT;
  wire fifo182_READ_OUTPUT;
  wire fifo183_READ_OUTPUT;
  wire fifo184_READ_OUTPUT;
  wire fifo185_READ_OUTPUT;
  wire fifo186_READ_OUTPUT;
  wire fifo187_READ_OUTPUT;
  wire fifo188_READ_OUTPUT;
  wire fifo189_READ_OUTPUT;
  wire fifo190_READ_OUTPUT;
  wire fifo191_READ_OUTPUT;
  wire fifo192_READ_OUTPUT;
  wire fifo193_READ_OUTPUT;
  wire fifo194_READ_OUTPUT;
  wire fifo195_READ_OUTPUT;
  wire fifo196_READ_OUTPUT;
  wire fifo197_READ_OUTPUT;
  wire fifo198_READ_OUTPUT;
  wire fifo199_READ_OUTPUT;
  wire fifo200_READ_OUTPUT;
  wire fifo201_READ_OUTPUT;
  wire fifo202_READ_OUTPUT;
  wire fifo203_READ_OUTPUT;
  wire fifo204_READ_OUTPUT;
  wire fifo205_READ_OUTPUT;
  wire fifo206_READ_OUTPUT;
  wire fifo207_READ_OUTPUT;
  wire fifo208_READ_OUTPUT;
  wire fifo209_READ_OUTPUT;
  wire fifo210_READ_OUTPUT;
  wire fifo211_READ_OUTPUT;
  wire fifo212_READ_OUTPUT;
  wire fifo213_READ_OUTPUT;
  wire fifo214_READ_OUTPUT;
  wire fifo215_READ_OUTPUT;
  wire fifo216_READ_OUTPUT;
  wire fifo217_READ_OUTPUT;
  wire fifo218_READ_OUTPUT;
  wire fifo219_READ_OUTPUT;
  wire fifo220_READ_OUTPUT;
  wire fifo221_READ_OUTPUT;
  wire fifo222_READ_OUTPUT;
  wire fifo223_READ_OUTPUT;
  wire fifo224_READ_OUTPUT;
  wire fifo225_READ_OUTPUT;
  wire fifo226_READ_OUTPUT;
  wire fifo227_READ_OUTPUT;
  wire fifo228_READ_OUTPUT;
  wire fifo229_READ_OUTPUT;
  wire fifo230_READ_OUTPUT;
  wire fifo231_READ_OUTPUT;
  wire fifo232_READ_OUTPUT;
  wire fifo233_READ_OUTPUT;
  wire fifo234_READ_OUTPUT;
  wire fifo235_READ_OUTPUT;
  wire fifo236_READ_OUTPUT;
  wire fifo237_READ_OUTPUT;
  wire fifo238_READ_OUTPUT;
  wire fifo239_READ_OUTPUT;
  wire fifo240_READ_OUTPUT;
  wire fifo241_READ_OUTPUT;
  wire fifo242_READ_OUTPUT;
  wire fifo243_READ_OUTPUT;
  wire fifo244_READ_OUTPUT;
  wire fifo245_READ_OUTPUT;
  wire fifo246_READ_OUTPUT;
  wire fifo247_READ_OUTPUT;
  wire fifo248_READ_OUTPUT;
  wire fifo249_READ_OUTPUT;
  wire fifo250_READ_OUTPUT;
  wire fifo251_READ_OUTPUT;
  wire fifo252_READ_OUTPUT;
  wire fifo253_READ_OUTPUT;
  wire fifo254_READ_OUTPUT;
  wire fifo255_READ_OUTPUT;
  wire fifo256_READ_OUTPUT;
  wire [7:0] writeAddr_GET_OUTPUT;
  wire unnamedunary6699USEDMULTIPLEunary = {(~{(writeAddr_GET_OUTPUT==readAddr_GET_OUTPUT)})};
  always @(posedge CLK) begin if(unnamedunary6699USEDMULTIPLEunary == 1'b0 && popFront_valid==1'b1 && CE_pop==1'b1) begin $display("%s: attempting to pop from an empty fifo",INSTANCE_NAME);$finish();  end end
  wire [7:0] readAddr_SETBY_OUTPUT;
  assign popFront = {fifo256_READ_OUTPUT,fifo255_READ_OUTPUT,fifo254_READ_OUTPUT,fifo253_READ_OUTPUT,fifo252_READ_OUTPUT,fifo251_READ_OUTPUT,fifo250_READ_OUTPUT,fifo249_READ_OUTPUT,fifo248_READ_OUTPUT,fifo247_READ_OUTPUT,fifo246_READ_OUTPUT,fifo245_READ_OUTPUT,fifo244_READ_OUTPUT,fifo243_READ_OUTPUT,fifo242_READ_OUTPUT,fifo241_READ_OUTPUT,fifo240_READ_OUTPUT,fifo239_READ_OUTPUT,fifo238_READ_OUTPUT,fifo237_READ_OUTPUT,fifo236_READ_OUTPUT,fifo235_READ_OUTPUT,fifo234_READ_OUTPUT,fifo233_READ_OUTPUT,fifo232_READ_OUTPUT,fifo231_READ_OUTPUT,fifo230_READ_OUTPUT,fifo229_READ_OUTPUT,fifo228_READ_OUTPUT,fifo227_READ_OUTPUT,fifo226_READ_OUTPUT,fifo225_READ_OUTPUT,fifo224_READ_OUTPUT,fifo223_READ_OUTPUT,fifo222_READ_OUTPUT,fifo221_READ_OUTPUT,fifo220_READ_OUTPUT,fifo219_READ_OUTPUT,fifo218_READ_OUTPUT,fifo217_READ_OUTPUT,fifo216_READ_OUTPUT,fifo215_READ_OUTPUT,fifo214_READ_OUTPUT,fifo213_READ_OUTPUT,fifo212_READ_OUTPUT,fifo211_READ_OUTPUT,fifo210_READ_OUTPUT,fifo209_READ_OUTPUT,fifo208_READ_OUTPUT,fifo207_READ_OUTPUT,fifo206_READ_OUTPUT,fifo205_READ_OUTPUT,fifo204_READ_OUTPUT,fifo203_READ_OUTPUT,fifo202_READ_OUTPUT,fifo201_READ_OUTPUT,fifo200_READ_OUTPUT,fifo199_READ_OUTPUT,fifo198_READ_OUTPUT,fifo197_READ_OUTPUT,fifo196_READ_OUTPUT,fifo195_READ_OUTPUT,fifo194_READ_OUTPUT,fifo193_READ_OUTPUT,fifo192_READ_OUTPUT,fifo191_READ_OUTPUT,fifo190_READ_OUTPUT,fifo189_READ_OUTPUT,fifo188_READ_OUTPUT,fifo187_READ_OUTPUT,fifo186_READ_OUTPUT,fifo185_READ_OUTPUT,fifo184_READ_OUTPUT,fifo183_READ_OUTPUT,fifo182_READ_OUTPUT,fifo181_READ_OUTPUT,fifo180_READ_OUTPUT,fifo179_READ_OUTPUT,fifo178_READ_OUTPUT,fifo177_READ_OUTPUT,fifo176_READ_OUTPUT,fifo175_READ_OUTPUT,fifo174_READ_OUTPUT,fifo173_READ_OUTPUT,fifo172_READ_OUTPUT,fifo171_READ_OUTPUT,fifo170_READ_OUTPUT,fifo169_READ_OUTPUT,fifo168_READ_OUTPUT,fifo167_READ_OUTPUT,fifo166_READ_OUTPUT,fifo165_READ_OUTPUT,fifo164_READ_OUTPUT,fifo163_READ_OUTPUT,fifo162_READ_OUTPUT,fifo161_READ_OUTPUT,fifo160_READ_OUTPUT,fifo159_READ_OUTPUT,fifo158_READ_OUTPUT,fifo157_READ_OUTPUT,fifo156_READ_OUTPUT,fifo155_READ_OUTPUT,fifo154_READ_OUTPUT,fifo153_READ_OUTPUT,fifo152_READ_OUTPUT,fifo151_READ_OUTPUT,fifo150_READ_OUTPUT,fifo149_READ_OUTPUT,fifo148_READ_OUTPUT,fifo147_READ_OUTPUT,fifo146_READ_OUTPUT,fifo145_READ_OUTPUT,fifo144_READ_OUTPUT,fifo143_READ_OUTPUT,fifo142_READ_OUTPUT,fifo141_READ_OUTPUT,fifo140_READ_OUTPUT,fifo139_READ_OUTPUT,fifo138_READ_OUTPUT,fifo137_READ_OUTPUT,fifo136_READ_OUTPUT,fifo135_READ_OUTPUT,fifo134_READ_OUTPUT,fifo133_READ_OUTPUT,fifo132_READ_OUTPUT,fifo131_READ_OUTPUT,fifo130_READ_OUTPUT,fifo129_READ_OUTPUT,fifo128_READ_OUTPUT,fifo127_READ_OUTPUT,fifo126_READ_OUTPUT,fifo125_READ_OUTPUT,fifo124_READ_OUTPUT,fifo123_READ_OUTPUT,fifo122_READ_OUTPUT,fifo121_READ_OUTPUT,fifo120_READ_OUTPUT,fifo119_READ_OUTPUT,fifo118_READ_OUTPUT,fifo117_READ_OUTPUT,fifo116_READ_OUTPUT,fifo115_READ_OUTPUT,fifo114_READ_OUTPUT,fifo113_READ_OUTPUT,fifo112_READ_OUTPUT,fifo111_READ_OUTPUT,fifo110_READ_OUTPUT,fifo109_READ_OUTPUT,fifo108_READ_OUTPUT,fifo107_READ_OUTPUT,fifo106_READ_OUTPUT,fifo105_READ_OUTPUT,fifo104_READ_OUTPUT,fifo103_READ_OUTPUT,fifo102_READ_OUTPUT,fifo101_READ_OUTPUT,fifo100_READ_OUTPUT,fifo99_READ_OUTPUT,fifo98_READ_OUTPUT,fifo97_READ_OUTPUT,fifo96_READ_OUTPUT,fifo95_READ_OUTPUT,fifo94_READ_OUTPUT,fifo93_READ_OUTPUT,fifo92_READ_OUTPUT,fifo91_READ_OUTPUT,fifo90_READ_OUTPUT,fifo89_READ_OUTPUT,fifo88_READ_OUTPUT,fifo87_READ_OUTPUT,fifo86_READ_OUTPUT,fifo85_READ_OUTPUT,fifo84_READ_OUTPUT,fifo83_READ_OUTPUT,fifo82_READ_OUTPUT,fifo81_READ_OUTPUT,fifo80_READ_OUTPUT,fifo79_READ_OUTPUT,fifo78_READ_OUTPUT,fifo77_READ_OUTPUT,fifo76_READ_OUTPUT,fifo75_READ_OUTPUT,fifo74_READ_OUTPUT,fifo73_READ_OUTPUT,fifo72_READ_OUTPUT,fifo71_READ_OUTPUT,fifo70_READ_OUTPUT,fifo69_READ_OUTPUT,fifo68_READ_OUTPUT,fifo67_READ_OUTPUT,fifo66_READ_OUTPUT,fifo65_READ_OUTPUT,fifo64_READ_OUTPUT,fifo63_READ_OUTPUT,fifo62_READ_OUTPUT,fifo61_READ_OUTPUT,fifo60_READ_OUTPUT,fifo59_READ_OUTPUT,fifo58_READ_OUTPUT,fifo57_READ_OUTPUT,fifo56_READ_OUTPUT,fifo55_READ_OUTPUT,fifo54_READ_OUTPUT,fifo53_READ_OUTPUT,fifo52_READ_OUTPUT,fifo51_READ_OUTPUT,fifo50_READ_OUTPUT,fifo49_READ_OUTPUT,fifo48_READ_OUTPUT,fifo47_READ_OUTPUT,fifo46_READ_OUTPUT,fifo45_READ_OUTPUT,fifo44_READ_OUTPUT,fifo43_READ_OUTPUT,fifo42_READ_OUTPUT,fifo41_READ_OUTPUT,fifo40_READ_OUTPUT,fifo39_READ_OUTPUT,fifo38_READ_OUTPUT,fifo37_READ_OUTPUT,fifo36_READ_OUTPUT,fifo35_READ_OUTPUT,fifo34_READ_OUTPUT,fifo33_READ_OUTPUT,fifo32_READ_OUTPUT,fifo31_READ_OUTPUT,fifo30_READ_OUTPUT,fifo29_READ_OUTPUT,fifo28_READ_OUTPUT,fifo27_READ_OUTPUT,fifo26_READ_OUTPUT,fifo25_READ_OUTPUT,fifo24_READ_OUTPUT,fifo23_READ_OUTPUT,fifo22_READ_OUTPUT,fifo21_READ_OUTPUT,fifo20_READ_OUTPUT,fifo19_READ_OUTPUT,fifo18_READ_OUTPUT,fifo17_READ_OUTPUT,fifo16_READ_OUTPUT,fifo15_READ_OUTPUT,fifo14_READ_OUTPUT,fifo13_READ_OUTPUT,fifo12_READ_OUTPUT,fifo11_READ_OUTPUT,fifo10_READ_OUTPUT,fifo9_READ_OUTPUT,fifo8_READ_OUTPUT,fifo7_READ_OUTPUT,fifo6_READ_OUTPUT,fifo5_READ_OUTPUT,fifo4_READ_OUTPUT,fifo3_READ_OUTPUT,fifo2_READ_OUTPUT,fifo1_READ_OUTPUT};
  wire [7:0] unnamedselect6690USEDMULTIPLEselect = (({((writeAddr_GET_OUTPUT)<(readAddr_GET_OUTPUT))})?({({((8'd128)-readAddr_GET_OUTPUT)}+writeAddr_GET_OUTPUT)}):({(writeAddr_GET_OUTPUT-readAddr_GET_OUTPUT)}));
  assign size = unnamedselect6690USEDMULTIPLEselect;
  reg readyReg;
    always @ (posedge CLK) begin readyReg <= {((unnamedselect6690USEDMULTIPLEselect)<((8'd125)))}; end
  assign ready = readyReg;
  always @(posedge CLK) begin if({((unnamedselect6690USEDMULTIPLEselect)<((8'd126)))} == 1'b0 && pushBack_valid==1'b1 && CE_push==1'b1) begin $display("%s: attempting to push to a full fifo",INSTANCE_NAME);$finish();  end end
  wire [7:0] writeAddr_SETBY_OUTPUT;
  wire [6:0] unnamedcast6707USEDMULTIPLEcast = writeAddr_GET_OUTPUT[6:0];
  assign hasData = unnamedunary6699USEDMULTIPLEunary;
  // function: popFront pure=false delay=0
  // function: size pure=true delay=0
  // function: pushBackReset pure=false delay=0
  // function: ready pure=true delay=0
  // function: pushBack pure=false delay=0
  // function: popFrontReset pure=false delay=0
  // function: hasData pure=true delay=0
  RegBy_incif_wrap127_incnil_CEtrue_initnil #(.INSTANCE_NAME("writeAddr")) writeAddr(.CLK(CLK), .set_valid(pushBackReset_valid), .CE(CE_push), .set_inp((8'd0)), .setby_valid(pushBack_valid), .setby_inp((1'd1)), .SETBY_OUTPUT(writeAddr_SETBY_OUTPUT), .GET_OUTPUT(writeAddr_GET_OUTPUT));
  RegBy_incif_wrap127_incnil_CEtrue_initnil #(.INSTANCE_NAME("readAddr")) readAddr(.CLK(CLK), .set_valid(popFrontReset_valid), .CE(CE_pop), .set_inp((8'd0)), .setby_valid(popFront_valid), .setby_inp((1'd1)), .SETBY_OUTPUT(readAddr_SETBY_OUTPUT), .GET_OUTPUT(readAddr_GET_OUTPUT));
  wire [7:0] fifo1_writeInput = {pushBack_input[0:0],unnamedcast6707USEDMULTIPLEcast};
wire fifo1_writeOut;
RAM128X1D fifo1  (
  .WCLK(CLK),
  .D(fifo1_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo1_writeOut),
  .DPO(fifo1_READ_OUTPUT),
  .A(fifo1_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo2_writeInput = {pushBack_input[1:1],unnamedcast6707USEDMULTIPLEcast};
wire fifo2_writeOut;
RAM128X1D fifo2  (
  .WCLK(CLK),
  .D(fifo2_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo2_writeOut),
  .DPO(fifo2_READ_OUTPUT),
  .A(fifo2_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo3_writeInput = {pushBack_input[2:2],unnamedcast6707USEDMULTIPLEcast};
wire fifo3_writeOut;
RAM128X1D fifo3  (
  .WCLK(CLK),
  .D(fifo3_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo3_writeOut),
  .DPO(fifo3_READ_OUTPUT),
  .A(fifo3_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo4_writeInput = {pushBack_input[3:3],unnamedcast6707USEDMULTIPLEcast};
wire fifo4_writeOut;
RAM128X1D fifo4  (
  .WCLK(CLK),
  .D(fifo4_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo4_writeOut),
  .DPO(fifo4_READ_OUTPUT),
  .A(fifo4_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo5_writeInput = {pushBack_input[4:4],unnamedcast6707USEDMULTIPLEcast};
wire fifo5_writeOut;
RAM128X1D fifo5  (
  .WCLK(CLK),
  .D(fifo5_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo5_writeOut),
  .DPO(fifo5_READ_OUTPUT),
  .A(fifo5_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo6_writeInput = {pushBack_input[5:5],unnamedcast6707USEDMULTIPLEcast};
wire fifo6_writeOut;
RAM128X1D fifo6  (
  .WCLK(CLK),
  .D(fifo6_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo6_writeOut),
  .DPO(fifo6_READ_OUTPUT),
  .A(fifo6_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo7_writeInput = {pushBack_input[6:6],unnamedcast6707USEDMULTIPLEcast};
wire fifo7_writeOut;
RAM128X1D fifo7  (
  .WCLK(CLK),
  .D(fifo7_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo7_writeOut),
  .DPO(fifo7_READ_OUTPUT),
  .A(fifo7_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo8_writeInput = {pushBack_input[7:7],unnamedcast6707USEDMULTIPLEcast};
wire fifo8_writeOut;
RAM128X1D fifo8  (
  .WCLK(CLK),
  .D(fifo8_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo8_writeOut),
  .DPO(fifo8_READ_OUTPUT),
  .A(fifo8_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo9_writeInput = {pushBack_input[8:8],unnamedcast6707USEDMULTIPLEcast};
wire fifo9_writeOut;
RAM128X1D fifo9  (
  .WCLK(CLK),
  .D(fifo9_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo9_writeOut),
  .DPO(fifo9_READ_OUTPUT),
  .A(fifo9_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo10_writeInput = {pushBack_input[9:9],unnamedcast6707USEDMULTIPLEcast};
wire fifo10_writeOut;
RAM128X1D fifo10  (
  .WCLK(CLK),
  .D(fifo10_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo10_writeOut),
  .DPO(fifo10_READ_OUTPUT),
  .A(fifo10_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo11_writeInput = {pushBack_input[10:10],unnamedcast6707USEDMULTIPLEcast};
wire fifo11_writeOut;
RAM128X1D fifo11  (
  .WCLK(CLK),
  .D(fifo11_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo11_writeOut),
  .DPO(fifo11_READ_OUTPUT),
  .A(fifo11_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo12_writeInput = {pushBack_input[11:11],unnamedcast6707USEDMULTIPLEcast};
wire fifo12_writeOut;
RAM128X1D fifo12  (
  .WCLK(CLK),
  .D(fifo12_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo12_writeOut),
  .DPO(fifo12_READ_OUTPUT),
  .A(fifo12_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo13_writeInput = {pushBack_input[12:12],unnamedcast6707USEDMULTIPLEcast};
wire fifo13_writeOut;
RAM128X1D fifo13  (
  .WCLK(CLK),
  .D(fifo13_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo13_writeOut),
  .DPO(fifo13_READ_OUTPUT),
  .A(fifo13_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo14_writeInput = {pushBack_input[13:13],unnamedcast6707USEDMULTIPLEcast};
wire fifo14_writeOut;
RAM128X1D fifo14  (
  .WCLK(CLK),
  .D(fifo14_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo14_writeOut),
  .DPO(fifo14_READ_OUTPUT),
  .A(fifo14_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo15_writeInput = {pushBack_input[14:14],unnamedcast6707USEDMULTIPLEcast};
wire fifo15_writeOut;
RAM128X1D fifo15  (
  .WCLK(CLK),
  .D(fifo15_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo15_writeOut),
  .DPO(fifo15_READ_OUTPUT),
  .A(fifo15_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo16_writeInput = {pushBack_input[15:15],unnamedcast6707USEDMULTIPLEcast};
wire fifo16_writeOut;
RAM128X1D fifo16  (
  .WCLK(CLK),
  .D(fifo16_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo16_writeOut),
  .DPO(fifo16_READ_OUTPUT),
  .A(fifo16_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo17_writeInput = {pushBack_input[16:16],unnamedcast6707USEDMULTIPLEcast};
wire fifo17_writeOut;
RAM128X1D fifo17  (
  .WCLK(CLK),
  .D(fifo17_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo17_writeOut),
  .DPO(fifo17_READ_OUTPUT),
  .A(fifo17_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo18_writeInput = {pushBack_input[17:17],unnamedcast6707USEDMULTIPLEcast};
wire fifo18_writeOut;
RAM128X1D fifo18  (
  .WCLK(CLK),
  .D(fifo18_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo18_writeOut),
  .DPO(fifo18_READ_OUTPUT),
  .A(fifo18_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo19_writeInput = {pushBack_input[18:18],unnamedcast6707USEDMULTIPLEcast};
wire fifo19_writeOut;
RAM128X1D fifo19  (
  .WCLK(CLK),
  .D(fifo19_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo19_writeOut),
  .DPO(fifo19_READ_OUTPUT),
  .A(fifo19_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo20_writeInput = {pushBack_input[19:19],unnamedcast6707USEDMULTIPLEcast};
wire fifo20_writeOut;
RAM128X1D fifo20  (
  .WCLK(CLK),
  .D(fifo20_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo20_writeOut),
  .DPO(fifo20_READ_OUTPUT),
  .A(fifo20_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo21_writeInput = {pushBack_input[20:20],unnamedcast6707USEDMULTIPLEcast};
wire fifo21_writeOut;
RAM128X1D fifo21  (
  .WCLK(CLK),
  .D(fifo21_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo21_writeOut),
  .DPO(fifo21_READ_OUTPUT),
  .A(fifo21_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo22_writeInput = {pushBack_input[21:21],unnamedcast6707USEDMULTIPLEcast};
wire fifo22_writeOut;
RAM128X1D fifo22  (
  .WCLK(CLK),
  .D(fifo22_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo22_writeOut),
  .DPO(fifo22_READ_OUTPUT),
  .A(fifo22_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo23_writeInput = {pushBack_input[22:22],unnamedcast6707USEDMULTIPLEcast};
wire fifo23_writeOut;
RAM128X1D fifo23  (
  .WCLK(CLK),
  .D(fifo23_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo23_writeOut),
  .DPO(fifo23_READ_OUTPUT),
  .A(fifo23_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo24_writeInput = {pushBack_input[23:23],unnamedcast6707USEDMULTIPLEcast};
wire fifo24_writeOut;
RAM128X1D fifo24  (
  .WCLK(CLK),
  .D(fifo24_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo24_writeOut),
  .DPO(fifo24_READ_OUTPUT),
  .A(fifo24_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo25_writeInput = {pushBack_input[24:24],unnamedcast6707USEDMULTIPLEcast};
wire fifo25_writeOut;
RAM128X1D fifo25  (
  .WCLK(CLK),
  .D(fifo25_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo25_writeOut),
  .DPO(fifo25_READ_OUTPUT),
  .A(fifo25_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo26_writeInput = {pushBack_input[25:25],unnamedcast6707USEDMULTIPLEcast};
wire fifo26_writeOut;
RAM128X1D fifo26  (
  .WCLK(CLK),
  .D(fifo26_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo26_writeOut),
  .DPO(fifo26_READ_OUTPUT),
  .A(fifo26_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo27_writeInput = {pushBack_input[26:26],unnamedcast6707USEDMULTIPLEcast};
wire fifo27_writeOut;
RAM128X1D fifo27  (
  .WCLK(CLK),
  .D(fifo27_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo27_writeOut),
  .DPO(fifo27_READ_OUTPUT),
  .A(fifo27_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo28_writeInput = {pushBack_input[27:27],unnamedcast6707USEDMULTIPLEcast};
wire fifo28_writeOut;
RAM128X1D fifo28  (
  .WCLK(CLK),
  .D(fifo28_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo28_writeOut),
  .DPO(fifo28_READ_OUTPUT),
  .A(fifo28_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo29_writeInput = {pushBack_input[28:28],unnamedcast6707USEDMULTIPLEcast};
wire fifo29_writeOut;
RAM128X1D fifo29  (
  .WCLK(CLK),
  .D(fifo29_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo29_writeOut),
  .DPO(fifo29_READ_OUTPUT),
  .A(fifo29_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo30_writeInput = {pushBack_input[29:29],unnamedcast6707USEDMULTIPLEcast};
wire fifo30_writeOut;
RAM128X1D fifo30  (
  .WCLK(CLK),
  .D(fifo30_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo30_writeOut),
  .DPO(fifo30_READ_OUTPUT),
  .A(fifo30_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo31_writeInput = {pushBack_input[30:30],unnamedcast6707USEDMULTIPLEcast};
wire fifo31_writeOut;
RAM128X1D fifo31  (
  .WCLK(CLK),
  .D(fifo31_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo31_writeOut),
  .DPO(fifo31_READ_OUTPUT),
  .A(fifo31_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo32_writeInput = {pushBack_input[31:31],unnamedcast6707USEDMULTIPLEcast};
wire fifo32_writeOut;
RAM128X1D fifo32  (
  .WCLK(CLK),
  .D(fifo32_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo32_writeOut),
  .DPO(fifo32_READ_OUTPUT),
  .A(fifo32_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo33_writeInput = {pushBack_input[32:32],unnamedcast6707USEDMULTIPLEcast};
wire fifo33_writeOut;
RAM128X1D fifo33  (
  .WCLK(CLK),
  .D(fifo33_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo33_writeOut),
  .DPO(fifo33_READ_OUTPUT),
  .A(fifo33_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo34_writeInput = {pushBack_input[33:33],unnamedcast6707USEDMULTIPLEcast};
wire fifo34_writeOut;
RAM128X1D fifo34  (
  .WCLK(CLK),
  .D(fifo34_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo34_writeOut),
  .DPO(fifo34_READ_OUTPUT),
  .A(fifo34_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo35_writeInput = {pushBack_input[34:34],unnamedcast6707USEDMULTIPLEcast};
wire fifo35_writeOut;
RAM128X1D fifo35  (
  .WCLK(CLK),
  .D(fifo35_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo35_writeOut),
  .DPO(fifo35_READ_OUTPUT),
  .A(fifo35_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo36_writeInput = {pushBack_input[35:35],unnamedcast6707USEDMULTIPLEcast};
wire fifo36_writeOut;
RAM128X1D fifo36  (
  .WCLK(CLK),
  .D(fifo36_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo36_writeOut),
  .DPO(fifo36_READ_OUTPUT),
  .A(fifo36_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo37_writeInput = {pushBack_input[36:36],unnamedcast6707USEDMULTIPLEcast};
wire fifo37_writeOut;
RAM128X1D fifo37  (
  .WCLK(CLK),
  .D(fifo37_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo37_writeOut),
  .DPO(fifo37_READ_OUTPUT),
  .A(fifo37_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo38_writeInput = {pushBack_input[37:37],unnamedcast6707USEDMULTIPLEcast};
wire fifo38_writeOut;
RAM128X1D fifo38  (
  .WCLK(CLK),
  .D(fifo38_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo38_writeOut),
  .DPO(fifo38_READ_OUTPUT),
  .A(fifo38_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo39_writeInput = {pushBack_input[38:38],unnamedcast6707USEDMULTIPLEcast};
wire fifo39_writeOut;
RAM128X1D fifo39  (
  .WCLK(CLK),
  .D(fifo39_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo39_writeOut),
  .DPO(fifo39_READ_OUTPUT),
  .A(fifo39_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo40_writeInput = {pushBack_input[39:39],unnamedcast6707USEDMULTIPLEcast};
wire fifo40_writeOut;
RAM128X1D fifo40  (
  .WCLK(CLK),
  .D(fifo40_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo40_writeOut),
  .DPO(fifo40_READ_OUTPUT),
  .A(fifo40_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo41_writeInput = {pushBack_input[40:40],unnamedcast6707USEDMULTIPLEcast};
wire fifo41_writeOut;
RAM128X1D fifo41  (
  .WCLK(CLK),
  .D(fifo41_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo41_writeOut),
  .DPO(fifo41_READ_OUTPUT),
  .A(fifo41_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo42_writeInput = {pushBack_input[41:41],unnamedcast6707USEDMULTIPLEcast};
wire fifo42_writeOut;
RAM128X1D fifo42  (
  .WCLK(CLK),
  .D(fifo42_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo42_writeOut),
  .DPO(fifo42_READ_OUTPUT),
  .A(fifo42_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo43_writeInput = {pushBack_input[42:42],unnamedcast6707USEDMULTIPLEcast};
wire fifo43_writeOut;
RAM128X1D fifo43  (
  .WCLK(CLK),
  .D(fifo43_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo43_writeOut),
  .DPO(fifo43_READ_OUTPUT),
  .A(fifo43_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo44_writeInput = {pushBack_input[43:43],unnamedcast6707USEDMULTIPLEcast};
wire fifo44_writeOut;
RAM128X1D fifo44  (
  .WCLK(CLK),
  .D(fifo44_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo44_writeOut),
  .DPO(fifo44_READ_OUTPUT),
  .A(fifo44_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo45_writeInput = {pushBack_input[44:44],unnamedcast6707USEDMULTIPLEcast};
wire fifo45_writeOut;
RAM128X1D fifo45  (
  .WCLK(CLK),
  .D(fifo45_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo45_writeOut),
  .DPO(fifo45_READ_OUTPUT),
  .A(fifo45_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo46_writeInput = {pushBack_input[45:45],unnamedcast6707USEDMULTIPLEcast};
wire fifo46_writeOut;
RAM128X1D fifo46  (
  .WCLK(CLK),
  .D(fifo46_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo46_writeOut),
  .DPO(fifo46_READ_OUTPUT),
  .A(fifo46_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo47_writeInput = {pushBack_input[46:46],unnamedcast6707USEDMULTIPLEcast};
wire fifo47_writeOut;
RAM128X1D fifo47  (
  .WCLK(CLK),
  .D(fifo47_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo47_writeOut),
  .DPO(fifo47_READ_OUTPUT),
  .A(fifo47_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo48_writeInput = {pushBack_input[47:47],unnamedcast6707USEDMULTIPLEcast};
wire fifo48_writeOut;
RAM128X1D fifo48  (
  .WCLK(CLK),
  .D(fifo48_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo48_writeOut),
  .DPO(fifo48_READ_OUTPUT),
  .A(fifo48_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo49_writeInput = {pushBack_input[48:48],unnamedcast6707USEDMULTIPLEcast};
wire fifo49_writeOut;
RAM128X1D fifo49  (
  .WCLK(CLK),
  .D(fifo49_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo49_writeOut),
  .DPO(fifo49_READ_OUTPUT),
  .A(fifo49_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo50_writeInput = {pushBack_input[49:49],unnamedcast6707USEDMULTIPLEcast};
wire fifo50_writeOut;
RAM128X1D fifo50  (
  .WCLK(CLK),
  .D(fifo50_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo50_writeOut),
  .DPO(fifo50_READ_OUTPUT),
  .A(fifo50_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo51_writeInput = {pushBack_input[50:50],unnamedcast6707USEDMULTIPLEcast};
wire fifo51_writeOut;
RAM128X1D fifo51  (
  .WCLK(CLK),
  .D(fifo51_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo51_writeOut),
  .DPO(fifo51_READ_OUTPUT),
  .A(fifo51_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo52_writeInput = {pushBack_input[51:51],unnamedcast6707USEDMULTIPLEcast};
wire fifo52_writeOut;
RAM128X1D fifo52  (
  .WCLK(CLK),
  .D(fifo52_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo52_writeOut),
  .DPO(fifo52_READ_OUTPUT),
  .A(fifo52_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo53_writeInput = {pushBack_input[52:52],unnamedcast6707USEDMULTIPLEcast};
wire fifo53_writeOut;
RAM128X1D fifo53  (
  .WCLK(CLK),
  .D(fifo53_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo53_writeOut),
  .DPO(fifo53_READ_OUTPUT),
  .A(fifo53_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo54_writeInput = {pushBack_input[53:53],unnamedcast6707USEDMULTIPLEcast};
wire fifo54_writeOut;
RAM128X1D fifo54  (
  .WCLK(CLK),
  .D(fifo54_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo54_writeOut),
  .DPO(fifo54_READ_OUTPUT),
  .A(fifo54_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo55_writeInput = {pushBack_input[54:54],unnamedcast6707USEDMULTIPLEcast};
wire fifo55_writeOut;
RAM128X1D fifo55  (
  .WCLK(CLK),
  .D(fifo55_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo55_writeOut),
  .DPO(fifo55_READ_OUTPUT),
  .A(fifo55_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo56_writeInput = {pushBack_input[55:55],unnamedcast6707USEDMULTIPLEcast};
wire fifo56_writeOut;
RAM128X1D fifo56  (
  .WCLK(CLK),
  .D(fifo56_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo56_writeOut),
  .DPO(fifo56_READ_OUTPUT),
  .A(fifo56_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo57_writeInput = {pushBack_input[56:56],unnamedcast6707USEDMULTIPLEcast};
wire fifo57_writeOut;
RAM128X1D fifo57  (
  .WCLK(CLK),
  .D(fifo57_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo57_writeOut),
  .DPO(fifo57_READ_OUTPUT),
  .A(fifo57_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo58_writeInput = {pushBack_input[57:57],unnamedcast6707USEDMULTIPLEcast};
wire fifo58_writeOut;
RAM128X1D fifo58  (
  .WCLK(CLK),
  .D(fifo58_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo58_writeOut),
  .DPO(fifo58_READ_OUTPUT),
  .A(fifo58_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo59_writeInput = {pushBack_input[58:58],unnamedcast6707USEDMULTIPLEcast};
wire fifo59_writeOut;
RAM128X1D fifo59  (
  .WCLK(CLK),
  .D(fifo59_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo59_writeOut),
  .DPO(fifo59_READ_OUTPUT),
  .A(fifo59_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo60_writeInput = {pushBack_input[59:59],unnamedcast6707USEDMULTIPLEcast};
wire fifo60_writeOut;
RAM128X1D fifo60  (
  .WCLK(CLK),
  .D(fifo60_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo60_writeOut),
  .DPO(fifo60_READ_OUTPUT),
  .A(fifo60_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo61_writeInput = {pushBack_input[60:60],unnamedcast6707USEDMULTIPLEcast};
wire fifo61_writeOut;
RAM128X1D fifo61  (
  .WCLK(CLK),
  .D(fifo61_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo61_writeOut),
  .DPO(fifo61_READ_OUTPUT),
  .A(fifo61_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo62_writeInput = {pushBack_input[61:61],unnamedcast6707USEDMULTIPLEcast};
wire fifo62_writeOut;
RAM128X1D fifo62  (
  .WCLK(CLK),
  .D(fifo62_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo62_writeOut),
  .DPO(fifo62_READ_OUTPUT),
  .A(fifo62_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo63_writeInput = {pushBack_input[62:62],unnamedcast6707USEDMULTIPLEcast};
wire fifo63_writeOut;
RAM128X1D fifo63  (
  .WCLK(CLK),
  .D(fifo63_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo63_writeOut),
  .DPO(fifo63_READ_OUTPUT),
  .A(fifo63_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo64_writeInput = {pushBack_input[63:63],unnamedcast6707USEDMULTIPLEcast};
wire fifo64_writeOut;
RAM128X1D fifo64  (
  .WCLK(CLK),
  .D(fifo64_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo64_writeOut),
  .DPO(fifo64_READ_OUTPUT),
  .A(fifo64_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo65_writeInput = {pushBack_input[64:64],unnamedcast6707USEDMULTIPLEcast};
wire fifo65_writeOut;
RAM128X1D fifo65  (
  .WCLK(CLK),
  .D(fifo65_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo65_writeOut),
  .DPO(fifo65_READ_OUTPUT),
  .A(fifo65_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo66_writeInput = {pushBack_input[65:65],unnamedcast6707USEDMULTIPLEcast};
wire fifo66_writeOut;
RAM128X1D fifo66  (
  .WCLK(CLK),
  .D(fifo66_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo66_writeOut),
  .DPO(fifo66_READ_OUTPUT),
  .A(fifo66_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo67_writeInput = {pushBack_input[66:66],unnamedcast6707USEDMULTIPLEcast};
wire fifo67_writeOut;
RAM128X1D fifo67  (
  .WCLK(CLK),
  .D(fifo67_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo67_writeOut),
  .DPO(fifo67_READ_OUTPUT),
  .A(fifo67_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo68_writeInput = {pushBack_input[67:67],unnamedcast6707USEDMULTIPLEcast};
wire fifo68_writeOut;
RAM128X1D fifo68  (
  .WCLK(CLK),
  .D(fifo68_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo68_writeOut),
  .DPO(fifo68_READ_OUTPUT),
  .A(fifo68_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo69_writeInput = {pushBack_input[68:68],unnamedcast6707USEDMULTIPLEcast};
wire fifo69_writeOut;
RAM128X1D fifo69  (
  .WCLK(CLK),
  .D(fifo69_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo69_writeOut),
  .DPO(fifo69_READ_OUTPUT),
  .A(fifo69_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo70_writeInput = {pushBack_input[69:69],unnamedcast6707USEDMULTIPLEcast};
wire fifo70_writeOut;
RAM128X1D fifo70  (
  .WCLK(CLK),
  .D(fifo70_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo70_writeOut),
  .DPO(fifo70_READ_OUTPUT),
  .A(fifo70_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo71_writeInput = {pushBack_input[70:70],unnamedcast6707USEDMULTIPLEcast};
wire fifo71_writeOut;
RAM128X1D fifo71  (
  .WCLK(CLK),
  .D(fifo71_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo71_writeOut),
  .DPO(fifo71_READ_OUTPUT),
  .A(fifo71_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo72_writeInput = {pushBack_input[71:71],unnamedcast6707USEDMULTIPLEcast};
wire fifo72_writeOut;
RAM128X1D fifo72  (
  .WCLK(CLK),
  .D(fifo72_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo72_writeOut),
  .DPO(fifo72_READ_OUTPUT),
  .A(fifo72_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo73_writeInput = {pushBack_input[72:72],unnamedcast6707USEDMULTIPLEcast};
wire fifo73_writeOut;
RAM128X1D fifo73  (
  .WCLK(CLK),
  .D(fifo73_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo73_writeOut),
  .DPO(fifo73_READ_OUTPUT),
  .A(fifo73_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo74_writeInput = {pushBack_input[73:73],unnamedcast6707USEDMULTIPLEcast};
wire fifo74_writeOut;
RAM128X1D fifo74  (
  .WCLK(CLK),
  .D(fifo74_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo74_writeOut),
  .DPO(fifo74_READ_OUTPUT),
  .A(fifo74_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo75_writeInput = {pushBack_input[74:74],unnamedcast6707USEDMULTIPLEcast};
wire fifo75_writeOut;
RAM128X1D fifo75  (
  .WCLK(CLK),
  .D(fifo75_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo75_writeOut),
  .DPO(fifo75_READ_OUTPUT),
  .A(fifo75_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo76_writeInput = {pushBack_input[75:75],unnamedcast6707USEDMULTIPLEcast};
wire fifo76_writeOut;
RAM128X1D fifo76  (
  .WCLK(CLK),
  .D(fifo76_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo76_writeOut),
  .DPO(fifo76_READ_OUTPUT),
  .A(fifo76_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo77_writeInput = {pushBack_input[76:76],unnamedcast6707USEDMULTIPLEcast};
wire fifo77_writeOut;
RAM128X1D fifo77  (
  .WCLK(CLK),
  .D(fifo77_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo77_writeOut),
  .DPO(fifo77_READ_OUTPUT),
  .A(fifo77_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo78_writeInput = {pushBack_input[77:77],unnamedcast6707USEDMULTIPLEcast};
wire fifo78_writeOut;
RAM128X1D fifo78  (
  .WCLK(CLK),
  .D(fifo78_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo78_writeOut),
  .DPO(fifo78_READ_OUTPUT),
  .A(fifo78_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo79_writeInput = {pushBack_input[78:78],unnamedcast6707USEDMULTIPLEcast};
wire fifo79_writeOut;
RAM128X1D fifo79  (
  .WCLK(CLK),
  .D(fifo79_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo79_writeOut),
  .DPO(fifo79_READ_OUTPUT),
  .A(fifo79_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo80_writeInput = {pushBack_input[79:79],unnamedcast6707USEDMULTIPLEcast};
wire fifo80_writeOut;
RAM128X1D fifo80  (
  .WCLK(CLK),
  .D(fifo80_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo80_writeOut),
  .DPO(fifo80_READ_OUTPUT),
  .A(fifo80_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo81_writeInput = {pushBack_input[80:80],unnamedcast6707USEDMULTIPLEcast};
wire fifo81_writeOut;
RAM128X1D fifo81  (
  .WCLK(CLK),
  .D(fifo81_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo81_writeOut),
  .DPO(fifo81_READ_OUTPUT),
  .A(fifo81_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo82_writeInput = {pushBack_input[81:81],unnamedcast6707USEDMULTIPLEcast};
wire fifo82_writeOut;
RAM128X1D fifo82  (
  .WCLK(CLK),
  .D(fifo82_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo82_writeOut),
  .DPO(fifo82_READ_OUTPUT),
  .A(fifo82_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo83_writeInput = {pushBack_input[82:82],unnamedcast6707USEDMULTIPLEcast};
wire fifo83_writeOut;
RAM128X1D fifo83  (
  .WCLK(CLK),
  .D(fifo83_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo83_writeOut),
  .DPO(fifo83_READ_OUTPUT),
  .A(fifo83_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo84_writeInput = {pushBack_input[83:83],unnamedcast6707USEDMULTIPLEcast};
wire fifo84_writeOut;
RAM128X1D fifo84  (
  .WCLK(CLK),
  .D(fifo84_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo84_writeOut),
  .DPO(fifo84_READ_OUTPUT),
  .A(fifo84_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo85_writeInput = {pushBack_input[84:84],unnamedcast6707USEDMULTIPLEcast};
wire fifo85_writeOut;
RAM128X1D fifo85  (
  .WCLK(CLK),
  .D(fifo85_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo85_writeOut),
  .DPO(fifo85_READ_OUTPUT),
  .A(fifo85_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo86_writeInput = {pushBack_input[85:85],unnamedcast6707USEDMULTIPLEcast};
wire fifo86_writeOut;
RAM128X1D fifo86  (
  .WCLK(CLK),
  .D(fifo86_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo86_writeOut),
  .DPO(fifo86_READ_OUTPUT),
  .A(fifo86_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo87_writeInput = {pushBack_input[86:86],unnamedcast6707USEDMULTIPLEcast};
wire fifo87_writeOut;
RAM128X1D fifo87  (
  .WCLK(CLK),
  .D(fifo87_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo87_writeOut),
  .DPO(fifo87_READ_OUTPUT),
  .A(fifo87_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo88_writeInput = {pushBack_input[87:87],unnamedcast6707USEDMULTIPLEcast};
wire fifo88_writeOut;
RAM128X1D fifo88  (
  .WCLK(CLK),
  .D(fifo88_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo88_writeOut),
  .DPO(fifo88_READ_OUTPUT),
  .A(fifo88_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo89_writeInput = {pushBack_input[88:88],unnamedcast6707USEDMULTIPLEcast};
wire fifo89_writeOut;
RAM128X1D fifo89  (
  .WCLK(CLK),
  .D(fifo89_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo89_writeOut),
  .DPO(fifo89_READ_OUTPUT),
  .A(fifo89_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo90_writeInput = {pushBack_input[89:89],unnamedcast6707USEDMULTIPLEcast};
wire fifo90_writeOut;
RAM128X1D fifo90  (
  .WCLK(CLK),
  .D(fifo90_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo90_writeOut),
  .DPO(fifo90_READ_OUTPUT),
  .A(fifo90_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo91_writeInput = {pushBack_input[90:90],unnamedcast6707USEDMULTIPLEcast};
wire fifo91_writeOut;
RAM128X1D fifo91  (
  .WCLK(CLK),
  .D(fifo91_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo91_writeOut),
  .DPO(fifo91_READ_OUTPUT),
  .A(fifo91_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo92_writeInput = {pushBack_input[91:91],unnamedcast6707USEDMULTIPLEcast};
wire fifo92_writeOut;
RAM128X1D fifo92  (
  .WCLK(CLK),
  .D(fifo92_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo92_writeOut),
  .DPO(fifo92_READ_OUTPUT),
  .A(fifo92_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo93_writeInput = {pushBack_input[92:92],unnamedcast6707USEDMULTIPLEcast};
wire fifo93_writeOut;
RAM128X1D fifo93  (
  .WCLK(CLK),
  .D(fifo93_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo93_writeOut),
  .DPO(fifo93_READ_OUTPUT),
  .A(fifo93_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo94_writeInput = {pushBack_input[93:93],unnamedcast6707USEDMULTIPLEcast};
wire fifo94_writeOut;
RAM128X1D fifo94  (
  .WCLK(CLK),
  .D(fifo94_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo94_writeOut),
  .DPO(fifo94_READ_OUTPUT),
  .A(fifo94_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo95_writeInput = {pushBack_input[94:94],unnamedcast6707USEDMULTIPLEcast};
wire fifo95_writeOut;
RAM128X1D fifo95  (
  .WCLK(CLK),
  .D(fifo95_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo95_writeOut),
  .DPO(fifo95_READ_OUTPUT),
  .A(fifo95_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo96_writeInput = {pushBack_input[95:95],unnamedcast6707USEDMULTIPLEcast};
wire fifo96_writeOut;
RAM128X1D fifo96  (
  .WCLK(CLK),
  .D(fifo96_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo96_writeOut),
  .DPO(fifo96_READ_OUTPUT),
  .A(fifo96_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo97_writeInput = {pushBack_input[96:96],unnamedcast6707USEDMULTIPLEcast};
wire fifo97_writeOut;
RAM128X1D fifo97  (
  .WCLK(CLK),
  .D(fifo97_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo97_writeOut),
  .DPO(fifo97_READ_OUTPUT),
  .A(fifo97_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo98_writeInput = {pushBack_input[97:97],unnamedcast6707USEDMULTIPLEcast};
wire fifo98_writeOut;
RAM128X1D fifo98  (
  .WCLK(CLK),
  .D(fifo98_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo98_writeOut),
  .DPO(fifo98_READ_OUTPUT),
  .A(fifo98_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo99_writeInput = {pushBack_input[98:98],unnamedcast6707USEDMULTIPLEcast};
wire fifo99_writeOut;
RAM128X1D fifo99  (
  .WCLK(CLK),
  .D(fifo99_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo99_writeOut),
  .DPO(fifo99_READ_OUTPUT),
  .A(fifo99_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo100_writeInput = {pushBack_input[99:99],unnamedcast6707USEDMULTIPLEcast};
wire fifo100_writeOut;
RAM128X1D fifo100  (
  .WCLK(CLK),
  .D(fifo100_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo100_writeOut),
  .DPO(fifo100_READ_OUTPUT),
  .A(fifo100_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo101_writeInput = {pushBack_input[100:100],unnamedcast6707USEDMULTIPLEcast};
wire fifo101_writeOut;
RAM128X1D fifo101  (
  .WCLK(CLK),
  .D(fifo101_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo101_writeOut),
  .DPO(fifo101_READ_OUTPUT),
  .A(fifo101_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo102_writeInput = {pushBack_input[101:101],unnamedcast6707USEDMULTIPLEcast};
wire fifo102_writeOut;
RAM128X1D fifo102  (
  .WCLK(CLK),
  .D(fifo102_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo102_writeOut),
  .DPO(fifo102_READ_OUTPUT),
  .A(fifo102_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo103_writeInput = {pushBack_input[102:102],unnamedcast6707USEDMULTIPLEcast};
wire fifo103_writeOut;
RAM128X1D fifo103  (
  .WCLK(CLK),
  .D(fifo103_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo103_writeOut),
  .DPO(fifo103_READ_OUTPUT),
  .A(fifo103_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo104_writeInput = {pushBack_input[103:103],unnamedcast6707USEDMULTIPLEcast};
wire fifo104_writeOut;
RAM128X1D fifo104  (
  .WCLK(CLK),
  .D(fifo104_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo104_writeOut),
  .DPO(fifo104_READ_OUTPUT),
  .A(fifo104_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo105_writeInput = {pushBack_input[104:104],unnamedcast6707USEDMULTIPLEcast};
wire fifo105_writeOut;
RAM128X1D fifo105  (
  .WCLK(CLK),
  .D(fifo105_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo105_writeOut),
  .DPO(fifo105_READ_OUTPUT),
  .A(fifo105_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo106_writeInput = {pushBack_input[105:105],unnamedcast6707USEDMULTIPLEcast};
wire fifo106_writeOut;
RAM128X1D fifo106  (
  .WCLK(CLK),
  .D(fifo106_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo106_writeOut),
  .DPO(fifo106_READ_OUTPUT),
  .A(fifo106_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo107_writeInput = {pushBack_input[106:106],unnamedcast6707USEDMULTIPLEcast};
wire fifo107_writeOut;
RAM128X1D fifo107  (
  .WCLK(CLK),
  .D(fifo107_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo107_writeOut),
  .DPO(fifo107_READ_OUTPUT),
  .A(fifo107_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo108_writeInput = {pushBack_input[107:107],unnamedcast6707USEDMULTIPLEcast};
wire fifo108_writeOut;
RAM128X1D fifo108  (
  .WCLK(CLK),
  .D(fifo108_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo108_writeOut),
  .DPO(fifo108_READ_OUTPUT),
  .A(fifo108_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo109_writeInput = {pushBack_input[108:108],unnamedcast6707USEDMULTIPLEcast};
wire fifo109_writeOut;
RAM128X1D fifo109  (
  .WCLK(CLK),
  .D(fifo109_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo109_writeOut),
  .DPO(fifo109_READ_OUTPUT),
  .A(fifo109_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo110_writeInput = {pushBack_input[109:109],unnamedcast6707USEDMULTIPLEcast};
wire fifo110_writeOut;
RAM128X1D fifo110  (
  .WCLK(CLK),
  .D(fifo110_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo110_writeOut),
  .DPO(fifo110_READ_OUTPUT),
  .A(fifo110_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo111_writeInput = {pushBack_input[110:110],unnamedcast6707USEDMULTIPLEcast};
wire fifo111_writeOut;
RAM128X1D fifo111  (
  .WCLK(CLK),
  .D(fifo111_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo111_writeOut),
  .DPO(fifo111_READ_OUTPUT),
  .A(fifo111_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo112_writeInput = {pushBack_input[111:111],unnamedcast6707USEDMULTIPLEcast};
wire fifo112_writeOut;
RAM128X1D fifo112  (
  .WCLK(CLK),
  .D(fifo112_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo112_writeOut),
  .DPO(fifo112_READ_OUTPUT),
  .A(fifo112_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo113_writeInput = {pushBack_input[112:112],unnamedcast6707USEDMULTIPLEcast};
wire fifo113_writeOut;
RAM128X1D fifo113  (
  .WCLK(CLK),
  .D(fifo113_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo113_writeOut),
  .DPO(fifo113_READ_OUTPUT),
  .A(fifo113_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo114_writeInput = {pushBack_input[113:113],unnamedcast6707USEDMULTIPLEcast};
wire fifo114_writeOut;
RAM128X1D fifo114  (
  .WCLK(CLK),
  .D(fifo114_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo114_writeOut),
  .DPO(fifo114_READ_OUTPUT),
  .A(fifo114_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo115_writeInput = {pushBack_input[114:114],unnamedcast6707USEDMULTIPLEcast};
wire fifo115_writeOut;
RAM128X1D fifo115  (
  .WCLK(CLK),
  .D(fifo115_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo115_writeOut),
  .DPO(fifo115_READ_OUTPUT),
  .A(fifo115_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo116_writeInput = {pushBack_input[115:115],unnamedcast6707USEDMULTIPLEcast};
wire fifo116_writeOut;
RAM128X1D fifo116  (
  .WCLK(CLK),
  .D(fifo116_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo116_writeOut),
  .DPO(fifo116_READ_OUTPUT),
  .A(fifo116_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo117_writeInput = {pushBack_input[116:116],unnamedcast6707USEDMULTIPLEcast};
wire fifo117_writeOut;
RAM128X1D fifo117  (
  .WCLK(CLK),
  .D(fifo117_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo117_writeOut),
  .DPO(fifo117_READ_OUTPUT),
  .A(fifo117_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo118_writeInput = {pushBack_input[117:117],unnamedcast6707USEDMULTIPLEcast};
wire fifo118_writeOut;
RAM128X1D fifo118  (
  .WCLK(CLK),
  .D(fifo118_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo118_writeOut),
  .DPO(fifo118_READ_OUTPUT),
  .A(fifo118_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo119_writeInput = {pushBack_input[118:118],unnamedcast6707USEDMULTIPLEcast};
wire fifo119_writeOut;
RAM128X1D fifo119  (
  .WCLK(CLK),
  .D(fifo119_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo119_writeOut),
  .DPO(fifo119_READ_OUTPUT),
  .A(fifo119_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo120_writeInput = {pushBack_input[119:119],unnamedcast6707USEDMULTIPLEcast};
wire fifo120_writeOut;
RAM128X1D fifo120  (
  .WCLK(CLK),
  .D(fifo120_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo120_writeOut),
  .DPO(fifo120_READ_OUTPUT),
  .A(fifo120_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo121_writeInput = {pushBack_input[120:120],unnamedcast6707USEDMULTIPLEcast};
wire fifo121_writeOut;
RAM128X1D fifo121  (
  .WCLK(CLK),
  .D(fifo121_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo121_writeOut),
  .DPO(fifo121_READ_OUTPUT),
  .A(fifo121_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo122_writeInput = {pushBack_input[121:121],unnamedcast6707USEDMULTIPLEcast};
wire fifo122_writeOut;
RAM128X1D fifo122  (
  .WCLK(CLK),
  .D(fifo122_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo122_writeOut),
  .DPO(fifo122_READ_OUTPUT),
  .A(fifo122_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo123_writeInput = {pushBack_input[122:122],unnamedcast6707USEDMULTIPLEcast};
wire fifo123_writeOut;
RAM128X1D fifo123  (
  .WCLK(CLK),
  .D(fifo123_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo123_writeOut),
  .DPO(fifo123_READ_OUTPUT),
  .A(fifo123_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo124_writeInput = {pushBack_input[123:123],unnamedcast6707USEDMULTIPLEcast};
wire fifo124_writeOut;
RAM128X1D fifo124  (
  .WCLK(CLK),
  .D(fifo124_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo124_writeOut),
  .DPO(fifo124_READ_OUTPUT),
  .A(fifo124_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo125_writeInput = {pushBack_input[124:124],unnamedcast6707USEDMULTIPLEcast};
wire fifo125_writeOut;
RAM128X1D fifo125  (
  .WCLK(CLK),
  .D(fifo125_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo125_writeOut),
  .DPO(fifo125_READ_OUTPUT),
  .A(fifo125_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo126_writeInput = {pushBack_input[125:125],unnamedcast6707USEDMULTIPLEcast};
wire fifo126_writeOut;
RAM128X1D fifo126  (
  .WCLK(CLK),
  .D(fifo126_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo126_writeOut),
  .DPO(fifo126_READ_OUTPUT),
  .A(fifo126_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo127_writeInput = {pushBack_input[126:126],unnamedcast6707USEDMULTIPLEcast};
wire fifo127_writeOut;
RAM128X1D fifo127  (
  .WCLK(CLK),
  .D(fifo127_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo127_writeOut),
  .DPO(fifo127_READ_OUTPUT),
  .A(fifo127_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo128_writeInput = {pushBack_input[127:127],unnamedcast6707USEDMULTIPLEcast};
wire fifo128_writeOut;
RAM128X1D fifo128  (
  .WCLK(CLK),
  .D(fifo128_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo128_writeOut),
  .DPO(fifo128_READ_OUTPUT),
  .A(fifo128_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo129_writeInput = {pushBack_input[128:128],unnamedcast6707USEDMULTIPLEcast};
wire fifo129_writeOut;
RAM128X1D fifo129  (
  .WCLK(CLK),
  .D(fifo129_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo129_writeOut),
  .DPO(fifo129_READ_OUTPUT),
  .A(fifo129_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo130_writeInput = {pushBack_input[129:129],unnamedcast6707USEDMULTIPLEcast};
wire fifo130_writeOut;
RAM128X1D fifo130  (
  .WCLK(CLK),
  .D(fifo130_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo130_writeOut),
  .DPO(fifo130_READ_OUTPUT),
  .A(fifo130_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo131_writeInput = {pushBack_input[130:130],unnamedcast6707USEDMULTIPLEcast};
wire fifo131_writeOut;
RAM128X1D fifo131  (
  .WCLK(CLK),
  .D(fifo131_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo131_writeOut),
  .DPO(fifo131_READ_OUTPUT),
  .A(fifo131_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo132_writeInput = {pushBack_input[131:131],unnamedcast6707USEDMULTIPLEcast};
wire fifo132_writeOut;
RAM128X1D fifo132  (
  .WCLK(CLK),
  .D(fifo132_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo132_writeOut),
  .DPO(fifo132_READ_OUTPUT),
  .A(fifo132_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo133_writeInput = {pushBack_input[132:132],unnamedcast6707USEDMULTIPLEcast};
wire fifo133_writeOut;
RAM128X1D fifo133  (
  .WCLK(CLK),
  .D(fifo133_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo133_writeOut),
  .DPO(fifo133_READ_OUTPUT),
  .A(fifo133_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo134_writeInput = {pushBack_input[133:133],unnamedcast6707USEDMULTIPLEcast};
wire fifo134_writeOut;
RAM128X1D fifo134  (
  .WCLK(CLK),
  .D(fifo134_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo134_writeOut),
  .DPO(fifo134_READ_OUTPUT),
  .A(fifo134_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo135_writeInput = {pushBack_input[134:134],unnamedcast6707USEDMULTIPLEcast};
wire fifo135_writeOut;
RAM128X1D fifo135  (
  .WCLK(CLK),
  .D(fifo135_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo135_writeOut),
  .DPO(fifo135_READ_OUTPUT),
  .A(fifo135_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo136_writeInput = {pushBack_input[135:135],unnamedcast6707USEDMULTIPLEcast};
wire fifo136_writeOut;
RAM128X1D fifo136  (
  .WCLK(CLK),
  .D(fifo136_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo136_writeOut),
  .DPO(fifo136_READ_OUTPUT),
  .A(fifo136_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo137_writeInput = {pushBack_input[136:136],unnamedcast6707USEDMULTIPLEcast};
wire fifo137_writeOut;
RAM128X1D fifo137  (
  .WCLK(CLK),
  .D(fifo137_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo137_writeOut),
  .DPO(fifo137_READ_OUTPUT),
  .A(fifo137_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo138_writeInput = {pushBack_input[137:137],unnamedcast6707USEDMULTIPLEcast};
wire fifo138_writeOut;
RAM128X1D fifo138  (
  .WCLK(CLK),
  .D(fifo138_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo138_writeOut),
  .DPO(fifo138_READ_OUTPUT),
  .A(fifo138_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo139_writeInput = {pushBack_input[138:138],unnamedcast6707USEDMULTIPLEcast};
wire fifo139_writeOut;
RAM128X1D fifo139  (
  .WCLK(CLK),
  .D(fifo139_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo139_writeOut),
  .DPO(fifo139_READ_OUTPUT),
  .A(fifo139_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo140_writeInput = {pushBack_input[139:139],unnamedcast6707USEDMULTIPLEcast};
wire fifo140_writeOut;
RAM128X1D fifo140  (
  .WCLK(CLK),
  .D(fifo140_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo140_writeOut),
  .DPO(fifo140_READ_OUTPUT),
  .A(fifo140_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo141_writeInput = {pushBack_input[140:140],unnamedcast6707USEDMULTIPLEcast};
wire fifo141_writeOut;
RAM128X1D fifo141  (
  .WCLK(CLK),
  .D(fifo141_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo141_writeOut),
  .DPO(fifo141_READ_OUTPUT),
  .A(fifo141_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo142_writeInput = {pushBack_input[141:141],unnamedcast6707USEDMULTIPLEcast};
wire fifo142_writeOut;
RAM128X1D fifo142  (
  .WCLK(CLK),
  .D(fifo142_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo142_writeOut),
  .DPO(fifo142_READ_OUTPUT),
  .A(fifo142_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo143_writeInput = {pushBack_input[142:142],unnamedcast6707USEDMULTIPLEcast};
wire fifo143_writeOut;
RAM128X1D fifo143  (
  .WCLK(CLK),
  .D(fifo143_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo143_writeOut),
  .DPO(fifo143_READ_OUTPUT),
  .A(fifo143_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo144_writeInput = {pushBack_input[143:143],unnamedcast6707USEDMULTIPLEcast};
wire fifo144_writeOut;
RAM128X1D fifo144  (
  .WCLK(CLK),
  .D(fifo144_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo144_writeOut),
  .DPO(fifo144_READ_OUTPUT),
  .A(fifo144_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo145_writeInput = {pushBack_input[144:144],unnamedcast6707USEDMULTIPLEcast};
wire fifo145_writeOut;
RAM128X1D fifo145  (
  .WCLK(CLK),
  .D(fifo145_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo145_writeOut),
  .DPO(fifo145_READ_OUTPUT),
  .A(fifo145_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo146_writeInput = {pushBack_input[145:145],unnamedcast6707USEDMULTIPLEcast};
wire fifo146_writeOut;
RAM128X1D fifo146  (
  .WCLK(CLK),
  .D(fifo146_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo146_writeOut),
  .DPO(fifo146_READ_OUTPUT),
  .A(fifo146_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo147_writeInput = {pushBack_input[146:146],unnamedcast6707USEDMULTIPLEcast};
wire fifo147_writeOut;
RAM128X1D fifo147  (
  .WCLK(CLK),
  .D(fifo147_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo147_writeOut),
  .DPO(fifo147_READ_OUTPUT),
  .A(fifo147_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo148_writeInput = {pushBack_input[147:147],unnamedcast6707USEDMULTIPLEcast};
wire fifo148_writeOut;
RAM128X1D fifo148  (
  .WCLK(CLK),
  .D(fifo148_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo148_writeOut),
  .DPO(fifo148_READ_OUTPUT),
  .A(fifo148_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo149_writeInput = {pushBack_input[148:148],unnamedcast6707USEDMULTIPLEcast};
wire fifo149_writeOut;
RAM128X1D fifo149  (
  .WCLK(CLK),
  .D(fifo149_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo149_writeOut),
  .DPO(fifo149_READ_OUTPUT),
  .A(fifo149_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo150_writeInput = {pushBack_input[149:149],unnamedcast6707USEDMULTIPLEcast};
wire fifo150_writeOut;
RAM128X1D fifo150  (
  .WCLK(CLK),
  .D(fifo150_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo150_writeOut),
  .DPO(fifo150_READ_OUTPUT),
  .A(fifo150_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo151_writeInput = {pushBack_input[150:150],unnamedcast6707USEDMULTIPLEcast};
wire fifo151_writeOut;
RAM128X1D fifo151  (
  .WCLK(CLK),
  .D(fifo151_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo151_writeOut),
  .DPO(fifo151_READ_OUTPUT),
  .A(fifo151_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo152_writeInput = {pushBack_input[151:151],unnamedcast6707USEDMULTIPLEcast};
wire fifo152_writeOut;
RAM128X1D fifo152  (
  .WCLK(CLK),
  .D(fifo152_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo152_writeOut),
  .DPO(fifo152_READ_OUTPUT),
  .A(fifo152_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo153_writeInput = {pushBack_input[152:152],unnamedcast6707USEDMULTIPLEcast};
wire fifo153_writeOut;
RAM128X1D fifo153  (
  .WCLK(CLK),
  .D(fifo153_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo153_writeOut),
  .DPO(fifo153_READ_OUTPUT),
  .A(fifo153_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo154_writeInput = {pushBack_input[153:153],unnamedcast6707USEDMULTIPLEcast};
wire fifo154_writeOut;
RAM128X1D fifo154  (
  .WCLK(CLK),
  .D(fifo154_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo154_writeOut),
  .DPO(fifo154_READ_OUTPUT),
  .A(fifo154_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo155_writeInput = {pushBack_input[154:154],unnamedcast6707USEDMULTIPLEcast};
wire fifo155_writeOut;
RAM128X1D fifo155  (
  .WCLK(CLK),
  .D(fifo155_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo155_writeOut),
  .DPO(fifo155_READ_OUTPUT),
  .A(fifo155_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo156_writeInput = {pushBack_input[155:155],unnamedcast6707USEDMULTIPLEcast};
wire fifo156_writeOut;
RAM128X1D fifo156  (
  .WCLK(CLK),
  .D(fifo156_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo156_writeOut),
  .DPO(fifo156_READ_OUTPUT),
  .A(fifo156_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo157_writeInput = {pushBack_input[156:156],unnamedcast6707USEDMULTIPLEcast};
wire fifo157_writeOut;
RAM128X1D fifo157  (
  .WCLK(CLK),
  .D(fifo157_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo157_writeOut),
  .DPO(fifo157_READ_OUTPUT),
  .A(fifo157_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo158_writeInput = {pushBack_input[157:157],unnamedcast6707USEDMULTIPLEcast};
wire fifo158_writeOut;
RAM128X1D fifo158  (
  .WCLK(CLK),
  .D(fifo158_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo158_writeOut),
  .DPO(fifo158_READ_OUTPUT),
  .A(fifo158_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo159_writeInput = {pushBack_input[158:158],unnamedcast6707USEDMULTIPLEcast};
wire fifo159_writeOut;
RAM128X1D fifo159  (
  .WCLK(CLK),
  .D(fifo159_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo159_writeOut),
  .DPO(fifo159_READ_OUTPUT),
  .A(fifo159_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo160_writeInput = {pushBack_input[159:159],unnamedcast6707USEDMULTIPLEcast};
wire fifo160_writeOut;
RAM128X1D fifo160  (
  .WCLK(CLK),
  .D(fifo160_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo160_writeOut),
  .DPO(fifo160_READ_OUTPUT),
  .A(fifo160_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo161_writeInput = {pushBack_input[160:160],unnamedcast6707USEDMULTIPLEcast};
wire fifo161_writeOut;
RAM128X1D fifo161  (
  .WCLK(CLK),
  .D(fifo161_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo161_writeOut),
  .DPO(fifo161_READ_OUTPUT),
  .A(fifo161_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo162_writeInput = {pushBack_input[161:161],unnamedcast6707USEDMULTIPLEcast};
wire fifo162_writeOut;
RAM128X1D fifo162  (
  .WCLK(CLK),
  .D(fifo162_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo162_writeOut),
  .DPO(fifo162_READ_OUTPUT),
  .A(fifo162_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo163_writeInput = {pushBack_input[162:162],unnamedcast6707USEDMULTIPLEcast};
wire fifo163_writeOut;
RAM128X1D fifo163  (
  .WCLK(CLK),
  .D(fifo163_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo163_writeOut),
  .DPO(fifo163_READ_OUTPUT),
  .A(fifo163_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo164_writeInput = {pushBack_input[163:163],unnamedcast6707USEDMULTIPLEcast};
wire fifo164_writeOut;
RAM128X1D fifo164  (
  .WCLK(CLK),
  .D(fifo164_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo164_writeOut),
  .DPO(fifo164_READ_OUTPUT),
  .A(fifo164_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo165_writeInput = {pushBack_input[164:164],unnamedcast6707USEDMULTIPLEcast};
wire fifo165_writeOut;
RAM128X1D fifo165  (
  .WCLK(CLK),
  .D(fifo165_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo165_writeOut),
  .DPO(fifo165_READ_OUTPUT),
  .A(fifo165_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo166_writeInput = {pushBack_input[165:165],unnamedcast6707USEDMULTIPLEcast};
wire fifo166_writeOut;
RAM128X1D fifo166  (
  .WCLK(CLK),
  .D(fifo166_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo166_writeOut),
  .DPO(fifo166_READ_OUTPUT),
  .A(fifo166_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo167_writeInput = {pushBack_input[166:166],unnamedcast6707USEDMULTIPLEcast};
wire fifo167_writeOut;
RAM128X1D fifo167  (
  .WCLK(CLK),
  .D(fifo167_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo167_writeOut),
  .DPO(fifo167_READ_OUTPUT),
  .A(fifo167_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo168_writeInput = {pushBack_input[167:167],unnamedcast6707USEDMULTIPLEcast};
wire fifo168_writeOut;
RAM128X1D fifo168  (
  .WCLK(CLK),
  .D(fifo168_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo168_writeOut),
  .DPO(fifo168_READ_OUTPUT),
  .A(fifo168_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo169_writeInput = {pushBack_input[168:168],unnamedcast6707USEDMULTIPLEcast};
wire fifo169_writeOut;
RAM128X1D fifo169  (
  .WCLK(CLK),
  .D(fifo169_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo169_writeOut),
  .DPO(fifo169_READ_OUTPUT),
  .A(fifo169_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo170_writeInput = {pushBack_input[169:169],unnamedcast6707USEDMULTIPLEcast};
wire fifo170_writeOut;
RAM128X1D fifo170  (
  .WCLK(CLK),
  .D(fifo170_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo170_writeOut),
  .DPO(fifo170_READ_OUTPUT),
  .A(fifo170_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo171_writeInput = {pushBack_input[170:170],unnamedcast6707USEDMULTIPLEcast};
wire fifo171_writeOut;
RAM128X1D fifo171  (
  .WCLK(CLK),
  .D(fifo171_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo171_writeOut),
  .DPO(fifo171_READ_OUTPUT),
  .A(fifo171_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo172_writeInput = {pushBack_input[171:171],unnamedcast6707USEDMULTIPLEcast};
wire fifo172_writeOut;
RAM128X1D fifo172  (
  .WCLK(CLK),
  .D(fifo172_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo172_writeOut),
  .DPO(fifo172_READ_OUTPUT),
  .A(fifo172_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo173_writeInput = {pushBack_input[172:172],unnamedcast6707USEDMULTIPLEcast};
wire fifo173_writeOut;
RAM128X1D fifo173  (
  .WCLK(CLK),
  .D(fifo173_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo173_writeOut),
  .DPO(fifo173_READ_OUTPUT),
  .A(fifo173_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo174_writeInput = {pushBack_input[173:173],unnamedcast6707USEDMULTIPLEcast};
wire fifo174_writeOut;
RAM128X1D fifo174  (
  .WCLK(CLK),
  .D(fifo174_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo174_writeOut),
  .DPO(fifo174_READ_OUTPUT),
  .A(fifo174_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo175_writeInput = {pushBack_input[174:174],unnamedcast6707USEDMULTIPLEcast};
wire fifo175_writeOut;
RAM128X1D fifo175  (
  .WCLK(CLK),
  .D(fifo175_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo175_writeOut),
  .DPO(fifo175_READ_OUTPUT),
  .A(fifo175_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo176_writeInput = {pushBack_input[175:175],unnamedcast6707USEDMULTIPLEcast};
wire fifo176_writeOut;
RAM128X1D fifo176  (
  .WCLK(CLK),
  .D(fifo176_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo176_writeOut),
  .DPO(fifo176_READ_OUTPUT),
  .A(fifo176_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo177_writeInput = {pushBack_input[176:176],unnamedcast6707USEDMULTIPLEcast};
wire fifo177_writeOut;
RAM128X1D fifo177  (
  .WCLK(CLK),
  .D(fifo177_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo177_writeOut),
  .DPO(fifo177_READ_OUTPUT),
  .A(fifo177_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo178_writeInput = {pushBack_input[177:177],unnamedcast6707USEDMULTIPLEcast};
wire fifo178_writeOut;
RAM128X1D fifo178  (
  .WCLK(CLK),
  .D(fifo178_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo178_writeOut),
  .DPO(fifo178_READ_OUTPUT),
  .A(fifo178_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo179_writeInput = {pushBack_input[178:178],unnamedcast6707USEDMULTIPLEcast};
wire fifo179_writeOut;
RAM128X1D fifo179  (
  .WCLK(CLK),
  .D(fifo179_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo179_writeOut),
  .DPO(fifo179_READ_OUTPUT),
  .A(fifo179_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo180_writeInput = {pushBack_input[179:179],unnamedcast6707USEDMULTIPLEcast};
wire fifo180_writeOut;
RAM128X1D fifo180  (
  .WCLK(CLK),
  .D(fifo180_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo180_writeOut),
  .DPO(fifo180_READ_OUTPUT),
  .A(fifo180_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo181_writeInput = {pushBack_input[180:180],unnamedcast6707USEDMULTIPLEcast};
wire fifo181_writeOut;
RAM128X1D fifo181  (
  .WCLK(CLK),
  .D(fifo181_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo181_writeOut),
  .DPO(fifo181_READ_OUTPUT),
  .A(fifo181_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo182_writeInput = {pushBack_input[181:181],unnamedcast6707USEDMULTIPLEcast};
wire fifo182_writeOut;
RAM128X1D fifo182  (
  .WCLK(CLK),
  .D(fifo182_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo182_writeOut),
  .DPO(fifo182_READ_OUTPUT),
  .A(fifo182_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo183_writeInput = {pushBack_input[182:182],unnamedcast6707USEDMULTIPLEcast};
wire fifo183_writeOut;
RAM128X1D fifo183  (
  .WCLK(CLK),
  .D(fifo183_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo183_writeOut),
  .DPO(fifo183_READ_OUTPUT),
  .A(fifo183_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo184_writeInput = {pushBack_input[183:183],unnamedcast6707USEDMULTIPLEcast};
wire fifo184_writeOut;
RAM128X1D fifo184  (
  .WCLK(CLK),
  .D(fifo184_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo184_writeOut),
  .DPO(fifo184_READ_OUTPUT),
  .A(fifo184_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo185_writeInput = {pushBack_input[184:184],unnamedcast6707USEDMULTIPLEcast};
wire fifo185_writeOut;
RAM128X1D fifo185  (
  .WCLK(CLK),
  .D(fifo185_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo185_writeOut),
  .DPO(fifo185_READ_OUTPUT),
  .A(fifo185_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo186_writeInput = {pushBack_input[185:185],unnamedcast6707USEDMULTIPLEcast};
wire fifo186_writeOut;
RAM128X1D fifo186  (
  .WCLK(CLK),
  .D(fifo186_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo186_writeOut),
  .DPO(fifo186_READ_OUTPUT),
  .A(fifo186_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo187_writeInput = {pushBack_input[186:186],unnamedcast6707USEDMULTIPLEcast};
wire fifo187_writeOut;
RAM128X1D fifo187  (
  .WCLK(CLK),
  .D(fifo187_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo187_writeOut),
  .DPO(fifo187_READ_OUTPUT),
  .A(fifo187_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo188_writeInput = {pushBack_input[187:187],unnamedcast6707USEDMULTIPLEcast};
wire fifo188_writeOut;
RAM128X1D fifo188  (
  .WCLK(CLK),
  .D(fifo188_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo188_writeOut),
  .DPO(fifo188_READ_OUTPUT),
  .A(fifo188_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo189_writeInput = {pushBack_input[188:188],unnamedcast6707USEDMULTIPLEcast};
wire fifo189_writeOut;
RAM128X1D fifo189  (
  .WCLK(CLK),
  .D(fifo189_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo189_writeOut),
  .DPO(fifo189_READ_OUTPUT),
  .A(fifo189_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo190_writeInput = {pushBack_input[189:189],unnamedcast6707USEDMULTIPLEcast};
wire fifo190_writeOut;
RAM128X1D fifo190  (
  .WCLK(CLK),
  .D(fifo190_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo190_writeOut),
  .DPO(fifo190_READ_OUTPUT),
  .A(fifo190_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo191_writeInput = {pushBack_input[190:190],unnamedcast6707USEDMULTIPLEcast};
wire fifo191_writeOut;
RAM128X1D fifo191  (
  .WCLK(CLK),
  .D(fifo191_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo191_writeOut),
  .DPO(fifo191_READ_OUTPUT),
  .A(fifo191_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo192_writeInput = {pushBack_input[191:191],unnamedcast6707USEDMULTIPLEcast};
wire fifo192_writeOut;
RAM128X1D fifo192  (
  .WCLK(CLK),
  .D(fifo192_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo192_writeOut),
  .DPO(fifo192_READ_OUTPUT),
  .A(fifo192_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo193_writeInput = {pushBack_input[192:192],unnamedcast6707USEDMULTIPLEcast};
wire fifo193_writeOut;
RAM128X1D fifo193  (
  .WCLK(CLK),
  .D(fifo193_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo193_writeOut),
  .DPO(fifo193_READ_OUTPUT),
  .A(fifo193_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo194_writeInput = {pushBack_input[193:193],unnamedcast6707USEDMULTIPLEcast};
wire fifo194_writeOut;
RAM128X1D fifo194  (
  .WCLK(CLK),
  .D(fifo194_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo194_writeOut),
  .DPO(fifo194_READ_OUTPUT),
  .A(fifo194_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo195_writeInput = {pushBack_input[194:194],unnamedcast6707USEDMULTIPLEcast};
wire fifo195_writeOut;
RAM128X1D fifo195  (
  .WCLK(CLK),
  .D(fifo195_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo195_writeOut),
  .DPO(fifo195_READ_OUTPUT),
  .A(fifo195_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo196_writeInput = {pushBack_input[195:195],unnamedcast6707USEDMULTIPLEcast};
wire fifo196_writeOut;
RAM128X1D fifo196  (
  .WCLK(CLK),
  .D(fifo196_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo196_writeOut),
  .DPO(fifo196_READ_OUTPUT),
  .A(fifo196_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo197_writeInput = {pushBack_input[196:196],unnamedcast6707USEDMULTIPLEcast};
wire fifo197_writeOut;
RAM128X1D fifo197  (
  .WCLK(CLK),
  .D(fifo197_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo197_writeOut),
  .DPO(fifo197_READ_OUTPUT),
  .A(fifo197_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo198_writeInput = {pushBack_input[197:197],unnamedcast6707USEDMULTIPLEcast};
wire fifo198_writeOut;
RAM128X1D fifo198  (
  .WCLK(CLK),
  .D(fifo198_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo198_writeOut),
  .DPO(fifo198_READ_OUTPUT),
  .A(fifo198_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo199_writeInput = {pushBack_input[198:198],unnamedcast6707USEDMULTIPLEcast};
wire fifo199_writeOut;
RAM128X1D fifo199  (
  .WCLK(CLK),
  .D(fifo199_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo199_writeOut),
  .DPO(fifo199_READ_OUTPUT),
  .A(fifo199_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo200_writeInput = {pushBack_input[199:199],unnamedcast6707USEDMULTIPLEcast};
wire fifo200_writeOut;
RAM128X1D fifo200  (
  .WCLK(CLK),
  .D(fifo200_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo200_writeOut),
  .DPO(fifo200_READ_OUTPUT),
  .A(fifo200_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo201_writeInput = {pushBack_input[200:200],unnamedcast6707USEDMULTIPLEcast};
wire fifo201_writeOut;
RAM128X1D fifo201  (
  .WCLK(CLK),
  .D(fifo201_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo201_writeOut),
  .DPO(fifo201_READ_OUTPUT),
  .A(fifo201_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo202_writeInput = {pushBack_input[201:201],unnamedcast6707USEDMULTIPLEcast};
wire fifo202_writeOut;
RAM128X1D fifo202  (
  .WCLK(CLK),
  .D(fifo202_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo202_writeOut),
  .DPO(fifo202_READ_OUTPUT),
  .A(fifo202_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo203_writeInput = {pushBack_input[202:202],unnamedcast6707USEDMULTIPLEcast};
wire fifo203_writeOut;
RAM128X1D fifo203  (
  .WCLK(CLK),
  .D(fifo203_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo203_writeOut),
  .DPO(fifo203_READ_OUTPUT),
  .A(fifo203_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo204_writeInput = {pushBack_input[203:203],unnamedcast6707USEDMULTIPLEcast};
wire fifo204_writeOut;
RAM128X1D fifo204  (
  .WCLK(CLK),
  .D(fifo204_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo204_writeOut),
  .DPO(fifo204_READ_OUTPUT),
  .A(fifo204_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo205_writeInput = {pushBack_input[204:204],unnamedcast6707USEDMULTIPLEcast};
wire fifo205_writeOut;
RAM128X1D fifo205  (
  .WCLK(CLK),
  .D(fifo205_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo205_writeOut),
  .DPO(fifo205_READ_OUTPUT),
  .A(fifo205_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo206_writeInput = {pushBack_input[205:205],unnamedcast6707USEDMULTIPLEcast};
wire fifo206_writeOut;
RAM128X1D fifo206  (
  .WCLK(CLK),
  .D(fifo206_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo206_writeOut),
  .DPO(fifo206_READ_OUTPUT),
  .A(fifo206_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo207_writeInput = {pushBack_input[206:206],unnamedcast6707USEDMULTIPLEcast};
wire fifo207_writeOut;
RAM128X1D fifo207  (
  .WCLK(CLK),
  .D(fifo207_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo207_writeOut),
  .DPO(fifo207_READ_OUTPUT),
  .A(fifo207_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo208_writeInput = {pushBack_input[207:207],unnamedcast6707USEDMULTIPLEcast};
wire fifo208_writeOut;
RAM128X1D fifo208  (
  .WCLK(CLK),
  .D(fifo208_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo208_writeOut),
  .DPO(fifo208_READ_OUTPUT),
  .A(fifo208_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo209_writeInput = {pushBack_input[208:208],unnamedcast6707USEDMULTIPLEcast};
wire fifo209_writeOut;
RAM128X1D fifo209  (
  .WCLK(CLK),
  .D(fifo209_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo209_writeOut),
  .DPO(fifo209_READ_OUTPUT),
  .A(fifo209_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo210_writeInput = {pushBack_input[209:209],unnamedcast6707USEDMULTIPLEcast};
wire fifo210_writeOut;
RAM128X1D fifo210  (
  .WCLK(CLK),
  .D(fifo210_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo210_writeOut),
  .DPO(fifo210_READ_OUTPUT),
  .A(fifo210_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo211_writeInput = {pushBack_input[210:210],unnamedcast6707USEDMULTIPLEcast};
wire fifo211_writeOut;
RAM128X1D fifo211  (
  .WCLK(CLK),
  .D(fifo211_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo211_writeOut),
  .DPO(fifo211_READ_OUTPUT),
  .A(fifo211_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo212_writeInput = {pushBack_input[211:211],unnamedcast6707USEDMULTIPLEcast};
wire fifo212_writeOut;
RAM128X1D fifo212  (
  .WCLK(CLK),
  .D(fifo212_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo212_writeOut),
  .DPO(fifo212_READ_OUTPUT),
  .A(fifo212_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo213_writeInput = {pushBack_input[212:212],unnamedcast6707USEDMULTIPLEcast};
wire fifo213_writeOut;
RAM128X1D fifo213  (
  .WCLK(CLK),
  .D(fifo213_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo213_writeOut),
  .DPO(fifo213_READ_OUTPUT),
  .A(fifo213_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo214_writeInput = {pushBack_input[213:213],unnamedcast6707USEDMULTIPLEcast};
wire fifo214_writeOut;
RAM128X1D fifo214  (
  .WCLK(CLK),
  .D(fifo214_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo214_writeOut),
  .DPO(fifo214_READ_OUTPUT),
  .A(fifo214_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo215_writeInput = {pushBack_input[214:214],unnamedcast6707USEDMULTIPLEcast};
wire fifo215_writeOut;
RAM128X1D fifo215  (
  .WCLK(CLK),
  .D(fifo215_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo215_writeOut),
  .DPO(fifo215_READ_OUTPUT),
  .A(fifo215_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo216_writeInput = {pushBack_input[215:215],unnamedcast6707USEDMULTIPLEcast};
wire fifo216_writeOut;
RAM128X1D fifo216  (
  .WCLK(CLK),
  .D(fifo216_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo216_writeOut),
  .DPO(fifo216_READ_OUTPUT),
  .A(fifo216_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo217_writeInput = {pushBack_input[216:216],unnamedcast6707USEDMULTIPLEcast};
wire fifo217_writeOut;
RAM128X1D fifo217  (
  .WCLK(CLK),
  .D(fifo217_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo217_writeOut),
  .DPO(fifo217_READ_OUTPUT),
  .A(fifo217_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo218_writeInput = {pushBack_input[217:217],unnamedcast6707USEDMULTIPLEcast};
wire fifo218_writeOut;
RAM128X1D fifo218  (
  .WCLK(CLK),
  .D(fifo218_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo218_writeOut),
  .DPO(fifo218_READ_OUTPUT),
  .A(fifo218_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo219_writeInput = {pushBack_input[218:218],unnamedcast6707USEDMULTIPLEcast};
wire fifo219_writeOut;
RAM128X1D fifo219  (
  .WCLK(CLK),
  .D(fifo219_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo219_writeOut),
  .DPO(fifo219_READ_OUTPUT),
  .A(fifo219_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo220_writeInput = {pushBack_input[219:219],unnamedcast6707USEDMULTIPLEcast};
wire fifo220_writeOut;
RAM128X1D fifo220  (
  .WCLK(CLK),
  .D(fifo220_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo220_writeOut),
  .DPO(fifo220_READ_OUTPUT),
  .A(fifo220_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo221_writeInput = {pushBack_input[220:220],unnamedcast6707USEDMULTIPLEcast};
wire fifo221_writeOut;
RAM128X1D fifo221  (
  .WCLK(CLK),
  .D(fifo221_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo221_writeOut),
  .DPO(fifo221_READ_OUTPUT),
  .A(fifo221_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo222_writeInput = {pushBack_input[221:221],unnamedcast6707USEDMULTIPLEcast};
wire fifo222_writeOut;
RAM128X1D fifo222  (
  .WCLK(CLK),
  .D(fifo222_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo222_writeOut),
  .DPO(fifo222_READ_OUTPUT),
  .A(fifo222_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo223_writeInput = {pushBack_input[222:222],unnamedcast6707USEDMULTIPLEcast};
wire fifo223_writeOut;
RAM128X1D fifo223  (
  .WCLK(CLK),
  .D(fifo223_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo223_writeOut),
  .DPO(fifo223_READ_OUTPUT),
  .A(fifo223_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo224_writeInput = {pushBack_input[223:223],unnamedcast6707USEDMULTIPLEcast};
wire fifo224_writeOut;
RAM128X1D fifo224  (
  .WCLK(CLK),
  .D(fifo224_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo224_writeOut),
  .DPO(fifo224_READ_OUTPUT),
  .A(fifo224_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo225_writeInput = {pushBack_input[224:224],unnamedcast6707USEDMULTIPLEcast};
wire fifo225_writeOut;
RAM128X1D fifo225  (
  .WCLK(CLK),
  .D(fifo225_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo225_writeOut),
  .DPO(fifo225_READ_OUTPUT),
  .A(fifo225_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo226_writeInput = {pushBack_input[225:225],unnamedcast6707USEDMULTIPLEcast};
wire fifo226_writeOut;
RAM128X1D fifo226  (
  .WCLK(CLK),
  .D(fifo226_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo226_writeOut),
  .DPO(fifo226_READ_OUTPUT),
  .A(fifo226_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo227_writeInput = {pushBack_input[226:226],unnamedcast6707USEDMULTIPLEcast};
wire fifo227_writeOut;
RAM128X1D fifo227  (
  .WCLK(CLK),
  .D(fifo227_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo227_writeOut),
  .DPO(fifo227_READ_OUTPUT),
  .A(fifo227_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo228_writeInput = {pushBack_input[227:227],unnamedcast6707USEDMULTIPLEcast};
wire fifo228_writeOut;
RAM128X1D fifo228  (
  .WCLK(CLK),
  .D(fifo228_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo228_writeOut),
  .DPO(fifo228_READ_OUTPUT),
  .A(fifo228_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo229_writeInput = {pushBack_input[228:228],unnamedcast6707USEDMULTIPLEcast};
wire fifo229_writeOut;
RAM128X1D fifo229  (
  .WCLK(CLK),
  .D(fifo229_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo229_writeOut),
  .DPO(fifo229_READ_OUTPUT),
  .A(fifo229_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo230_writeInput = {pushBack_input[229:229],unnamedcast6707USEDMULTIPLEcast};
wire fifo230_writeOut;
RAM128X1D fifo230  (
  .WCLK(CLK),
  .D(fifo230_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo230_writeOut),
  .DPO(fifo230_READ_OUTPUT),
  .A(fifo230_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo231_writeInput = {pushBack_input[230:230],unnamedcast6707USEDMULTIPLEcast};
wire fifo231_writeOut;
RAM128X1D fifo231  (
  .WCLK(CLK),
  .D(fifo231_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo231_writeOut),
  .DPO(fifo231_READ_OUTPUT),
  .A(fifo231_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo232_writeInput = {pushBack_input[231:231],unnamedcast6707USEDMULTIPLEcast};
wire fifo232_writeOut;
RAM128X1D fifo232  (
  .WCLK(CLK),
  .D(fifo232_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo232_writeOut),
  .DPO(fifo232_READ_OUTPUT),
  .A(fifo232_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo233_writeInput = {pushBack_input[232:232],unnamedcast6707USEDMULTIPLEcast};
wire fifo233_writeOut;
RAM128X1D fifo233  (
  .WCLK(CLK),
  .D(fifo233_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo233_writeOut),
  .DPO(fifo233_READ_OUTPUT),
  .A(fifo233_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo234_writeInput = {pushBack_input[233:233],unnamedcast6707USEDMULTIPLEcast};
wire fifo234_writeOut;
RAM128X1D fifo234  (
  .WCLK(CLK),
  .D(fifo234_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo234_writeOut),
  .DPO(fifo234_READ_OUTPUT),
  .A(fifo234_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo235_writeInput = {pushBack_input[234:234],unnamedcast6707USEDMULTIPLEcast};
wire fifo235_writeOut;
RAM128X1D fifo235  (
  .WCLK(CLK),
  .D(fifo235_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo235_writeOut),
  .DPO(fifo235_READ_OUTPUT),
  .A(fifo235_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo236_writeInput = {pushBack_input[235:235],unnamedcast6707USEDMULTIPLEcast};
wire fifo236_writeOut;
RAM128X1D fifo236  (
  .WCLK(CLK),
  .D(fifo236_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo236_writeOut),
  .DPO(fifo236_READ_OUTPUT),
  .A(fifo236_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo237_writeInput = {pushBack_input[236:236],unnamedcast6707USEDMULTIPLEcast};
wire fifo237_writeOut;
RAM128X1D fifo237  (
  .WCLK(CLK),
  .D(fifo237_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo237_writeOut),
  .DPO(fifo237_READ_OUTPUT),
  .A(fifo237_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo238_writeInput = {pushBack_input[237:237],unnamedcast6707USEDMULTIPLEcast};
wire fifo238_writeOut;
RAM128X1D fifo238  (
  .WCLK(CLK),
  .D(fifo238_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo238_writeOut),
  .DPO(fifo238_READ_OUTPUT),
  .A(fifo238_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo239_writeInput = {pushBack_input[238:238],unnamedcast6707USEDMULTIPLEcast};
wire fifo239_writeOut;
RAM128X1D fifo239  (
  .WCLK(CLK),
  .D(fifo239_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo239_writeOut),
  .DPO(fifo239_READ_OUTPUT),
  .A(fifo239_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo240_writeInput = {pushBack_input[239:239],unnamedcast6707USEDMULTIPLEcast};
wire fifo240_writeOut;
RAM128X1D fifo240  (
  .WCLK(CLK),
  .D(fifo240_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo240_writeOut),
  .DPO(fifo240_READ_OUTPUT),
  .A(fifo240_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo241_writeInput = {pushBack_input[240:240],unnamedcast6707USEDMULTIPLEcast};
wire fifo241_writeOut;
RAM128X1D fifo241  (
  .WCLK(CLK),
  .D(fifo241_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo241_writeOut),
  .DPO(fifo241_READ_OUTPUT),
  .A(fifo241_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo242_writeInput = {pushBack_input[241:241],unnamedcast6707USEDMULTIPLEcast};
wire fifo242_writeOut;
RAM128X1D fifo242  (
  .WCLK(CLK),
  .D(fifo242_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo242_writeOut),
  .DPO(fifo242_READ_OUTPUT),
  .A(fifo242_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo243_writeInput = {pushBack_input[242:242],unnamedcast6707USEDMULTIPLEcast};
wire fifo243_writeOut;
RAM128X1D fifo243  (
  .WCLK(CLK),
  .D(fifo243_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo243_writeOut),
  .DPO(fifo243_READ_OUTPUT),
  .A(fifo243_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo244_writeInput = {pushBack_input[243:243],unnamedcast6707USEDMULTIPLEcast};
wire fifo244_writeOut;
RAM128X1D fifo244  (
  .WCLK(CLK),
  .D(fifo244_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo244_writeOut),
  .DPO(fifo244_READ_OUTPUT),
  .A(fifo244_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo245_writeInput = {pushBack_input[244:244],unnamedcast6707USEDMULTIPLEcast};
wire fifo245_writeOut;
RAM128X1D fifo245  (
  .WCLK(CLK),
  .D(fifo245_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo245_writeOut),
  .DPO(fifo245_READ_OUTPUT),
  .A(fifo245_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo246_writeInput = {pushBack_input[245:245],unnamedcast6707USEDMULTIPLEcast};
wire fifo246_writeOut;
RAM128X1D fifo246  (
  .WCLK(CLK),
  .D(fifo246_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo246_writeOut),
  .DPO(fifo246_READ_OUTPUT),
  .A(fifo246_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo247_writeInput = {pushBack_input[246:246],unnamedcast6707USEDMULTIPLEcast};
wire fifo247_writeOut;
RAM128X1D fifo247  (
  .WCLK(CLK),
  .D(fifo247_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo247_writeOut),
  .DPO(fifo247_READ_OUTPUT),
  .A(fifo247_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo248_writeInput = {pushBack_input[247:247],unnamedcast6707USEDMULTIPLEcast};
wire fifo248_writeOut;
RAM128X1D fifo248  (
  .WCLK(CLK),
  .D(fifo248_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo248_writeOut),
  .DPO(fifo248_READ_OUTPUT),
  .A(fifo248_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo249_writeInput = {pushBack_input[248:248],unnamedcast6707USEDMULTIPLEcast};
wire fifo249_writeOut;
RAM128X1D fifo249  (
  .WCLK(CLK),
  .D(fifo249_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo249_writeOut),
  .DPO(fifo249_READ_OUTPUT),
  .A(fifo249_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo250_writeInput = {pushBack_input[249:249],unnamedcast6707USEDMULTIPLEcast};
wire fifo250_writeOut;
RAM128X1D fifo250  (
  .WCLK(CLK),
  .D(fifo250_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo250_writeOut),
  .DPO(fifo250_READ_OUTPUT),
  .A(fifo250_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo251_writeInput = {pushBack_input[250:250],unnamedcast6707USEDMULTIPLEcast};
wire fifo251_writeOut;
RAM128X1D fifo251  (
  .WCLK(CLK),
  .D(fifo251_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo251_writeOut),
  .DPO(fifo251_READ_OUTPUT),
  .A(fifo251_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo252_writeInput = {pushBack_input[251:251],unnamedcast6707USEDMULTIPLEcast};
wire fifo252_writeOut;
RAM128X1D fifo252  (
  .WCLK(CLK),
  .D(fifo252_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo252_writeOut),
  .DPO(fifo252_READ_OUTPUT),
  .A(fifo252_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo253_writeInput = {pushBack_input[252:252],unnamedcast6707USEDMULTIPLEcast};
wire fifo253_writeOut;
RAM128X1D fifo253  (
  .WCLK(CLK),
  .D(fifo253_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo253_writeOut),
  .DPO(fifo253_READ_OUTPUT),
  .A(fifo253_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo254_writeInput = {pushBack_input[253:253],unnamedcast6707USEDMULTIPLEcast};
wire fifo254_writeOut;
RAM128X1D fifo254  (
  .WCLK(CLK),
  .D(fifo254_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo254_writeOut),
  .DPO(fifo254_READ_OUTPUT),
  .A(fifo254_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo255_writeInput = {pushBack_input[254:254],unnamedcast6707USEDMULTIPLEcast};
wire fifo255_writeOut;
RAM128X1D fifo255  (
  .WCLK(CLK),
  .D(fifo255_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo255_writeOut),
  .DPO(fifo255_READ_OUTPUT),
  .A(fifo255_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

  wire [7:0] fifo256_writeInput = {pushBack_input[255:255],unnamedcast6707USEDMULTIPLEcast};
wire fifo256_writeOut;
RAM128X1D fifo256  (
  .WCLK(CLK),
  .D(fifo256_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo256_writeOut),
  .DPO(fifo256_READ_OUTPUT),
  .A(fifo256_writeInput[6:0]),
  .DPRA(unnamedcast7992USEDMULTIPLEcast));

endmodule

module fifo_128_uint8_4_1__8_1_(input CLK, input load_valid, input load_CE, output [256:0] load_output, input store_reset_valid, input store_CE, output store_ready, input load_reset_valid, input store_valid, input [255:0] store_input);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(load_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_reset_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(load_reset_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store'", INSTANCE_NAME);  end end
  wire FIFO_hasData;
  wire [255:0] FIFO_popFront;
  assign load_output = {FIFO_hasData,FIFO_popFront};
  wire FIFO_ready;
  assign store_ready = FIFO_ready;
  // function: load pure=false delay=0
  // function: store_reset pure=false delay=0
  // function: store_ready pure=true delay=0
  // function: load_reset pure=false delay=0
  // function: store pure=false delay=0
  fifo_uint8_4_1__8_1_ #(.INSTANCE_NAME("FIFO")) FIFO(.CLK(CLK), .popFront_valid({(FIFO_hasData&&load_valid)}), .CE_pop(load_CE), .popFront(FIFO_popFront), .size(FIFO_size), .pushBackReset_valid(store_reset_valid), .CE_push(store_CE), .ready(FIFO_ready), .pushBack_valid(store_valid), .pushBack_input(store_input), .popFrontReset_valid(load_reset_valid), .hasData(FIFO_hasData));
endmodule

module LiftDecimate_fifo_128_uint8_4_1__8_1_(input CLK, input load_valid, input load_CE, input load_input, output [256:0] load_output, input store_reset_valid, input store_CE, output store_ready, output load_ready, input load_reset, input store_valid, input [255:0] store_input);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(load_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_reset_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(load_reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store'", INSTANCE_NAME);  end end
  wire unnamedcast11971USEDMULTIPLEcast = load_input;
  wire [256:0] LiftDecimate_inner_fifo_128_uint8_4_1__8_1__load_output;
  reg [255:0] unnamedcast11974_delay1_validunnamednull0_CEload_CE;  always @ (posedge CLK) begin if (load_CE) begin unnamedcast11974_delay1_validunnamednull0_CEload_CE <= (LiftDecimate_inner_fifo_128_uint8_4_1__8_1__load_output[255:0]); end end
  reg unnamedbinop11979_delay1_validunnamednull0_CEload_CE;  always @ (posedge CLK) begin if (load_CE) begin unnamedbinop11979_delay1_validunnamednull0_CEload_CE <= {((LiftDecimate_inner_fifo_128_uint8_4_1__8_1__load_output[256])&&unnamedcast11971USEDMULTIPLEcast)}; end end
  assign load_output = {unnamedbinop11979_delay1_validunnamednull0_CEload_CE,unnamedcast11974_delay1_validunnamednull0_CEload_CE};
  wire LiftDecimate_inner_fifo_128_uint8_4_1__8_1__store_ready;
  assign store_ready = LiftDecimate_inner_fifo_128_uint8_4_1__8_1__store_ready;
  assign load_ready = (1'd1);
  // function: load pure=false delay=1
  // function: store_reset pure=false delay=0
  // function: store_ready pure=true delay=0
  // function: load_ready pure=true delay=0
  // function: load_reset pure=false delay=0
  // function: store pure=false delay=0
  fifo_128_uint8_4_1__8_1_ #(.INSTANCE_NAME("LiftDecimate_inner_fifo_128_uint8_4_1__8_1_")) LiftDecimate_inner_fifo_128_uint8_4_1__8_1_(.CLK(CLK), .load_valid({(unnamedcast11971USEDMULTIPLEcast&&load_valid)}), .load_CE(load_CE), .load_output(LiftDecimate_inner_fifo_128_uint8_4_1__8_1__load_output), .store_reset_valid(store_reset_valid), .store_CE(store_CE), .store_ready(LiftDecimate_inner_fifo_128_uint8_4_1__8_1__store_ready), .load_reset_valid(load_reset), .store_valid(store_valid), .store_input(store_input));
endmodule

module RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1_(input CLK, input load_valid, input load_CE, input load_input, output [256:0] load_output, input store_reset, input CE, output store_ready, output load_ready, input load_reset, input store_valid, input [256:0] store_input, output store_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(load_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(load_reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store'", INSTANCE_NAME);  end end
  wire [256:0] RunIffReady_inner_load_output;
  assign load_output = RunIffReady_inner_load_output;
  wire RunIffReady_inner_store_ready;
  assign store_ready = RunIffReady_inner_store_ready;
  wire RunIffReady_inner_load_ready;
  assign load_ready = RunIffReady_inner_load_ready;
  wire unnamedbinop12050USEDMULTIPLEbinop = {({(RunIffReady_inner_store_ready&&(store_input[256]))}&&store_valid)};
  assign store_output = {unnamedbinop12050USEDMULTIPLEbinop};
  // function: load pure=false delay=1
  // function: store_reset pure=false delay=0
  // function: store_ready pure=true delay=0
  // function: load_ready pure=true delay=0
  // function: load_reset pure=false delay=0
  // function: store pure=false delay=0
  LiftDecimate_fifo_128_uint8_4_1__8_1_ #(.INSTANCE_NAME("RunIffReady_inner")) RunIffReady_inner(.CLK(CLK), .load_valid(load_valid), .load_CE(load_CE), .load_input(load_input), .load_output(RunIffReady_inner_load_output), .store_reset_valid(store_reset), .store_CE(CE), .store_ready(RunIffReady_inner_store_ready), .load_ready(RunIffReady_inner_load_ready), .load_reset(load_reset), .store_valid(unnamedbinop12050USEDMULTIPLEbinop), .store_input((store_input[255:0])));
endmodule

module LiftHandshake_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1_(input CLK, input load_input, output [256:0] load_output, input store_reset, input store_ready_downstream, output store_ready, input load_ready_downstream, output load_ready, input load_reset, input [256:0] store_input, output store_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire unnamedunary12087USEDMULTIPLEunary = {(~load_reset)};
  wire unnamedbinop12086USEDMULTIPLEbinop = {(load_reset||load_ready_downstream)};
  wire [256:0] inner_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1__load_output;
  wire load_validBitDelay_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1__pushPop_out;
  wire [256:0] unnamedtuple12097USEDMULTIPLEtuple = {{((inner_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1__load_output[256])&&load_validBitDelay_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1__pushPop_out)},(inner_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1__load_output[255:0])};
  always @(posedge CLK) begin if({(~{((unnamedtuple12097USEDMULTIPLEtuple[256])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: output valid bit should not be X!",INSTANCE_NAME); end end
  always @(posedge CLK) begin if({(~{(load_input===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign load_output = unnamedtuple12097USEDMULTIPLEtuple;
  wire unnamedbinop12115USEDMULTIPLEbinop = {(store_reset||store_ready_downstream)};
  wire inner_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1__store_ready;
  assign store_ready = {(inner_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1__store_ready&&store_ready_downstream)};
  wire inner_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1__load_ready;
  assign load_ready = {(inner_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1__load_ready&&load_ready_downstream)};
  wire unnamedunary12116USEDMULTIPLEunary = {(~store_reset)};
  wire [0:0] inner_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1__store_output;
  wire store_validBitDelay_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1__pushPop_out;
  wire [0:0] unnamedtuple12126USEDMULTIPLEtuple = {{(inner_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1__store_output&&store_validBitDelay_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1__pushPop_out)}};
  always @(posedge CLK) begin if({(~{(unnamedtuple12126USEDMULTIPLEtuple===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: output valid bit should not be X!",INSTANCE_NAME); end end
  always @(posedge CLK) begin if({(~{((store_input[256])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign store_output = unnamedtuple12126USEDMULTIPLEtuple;
  // function: load pure=false ONLY WIRE
  // function: store_reset pure=false ONLY WIRE
  // function: store_ready pure=true ONLY WIRE
  // function: load_ready pure=true ONLY WIRE
  // function: load_reset pure=false ONLY WIRE
  // function: store pure=false ONLY WIRE
  RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1_ #(.INSTANCE_NAME("inner_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1_")) inner_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1_(.CLK(CLK), .load_valid(unnamedunary12087USEDMULTIPLEunary), .load_CE(unnamedbinop12086USEDMULTIPLEbinop), .load_input(load_input), .load_output(inner_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1__load_output), .store_reset(store_reset), .CE(unnamedbinop12115USEDMULTIPLEbinop), .store_ready(inner_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1__store_ready), .load_ready(inner_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1__load_ready), .load_reset(load_reset), .store_valid(unnamedunary12116USEDMULTIPLEunary), .store_input(store_input), .store_output(inner_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1__store_output));
  ShiftRegister_1_CEtrue_TY1 #(.INSTANCE_NAME("load_validBitDelay_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1_")) load_validBitDelay_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1_(.CLK(CLK), .pushPop_valid(unnamedunary12087USEDMULTIPLEunary), .CE(unnamedbinop12086USEDMULTIPLEbinop), .sr_input((1'd1)), .pushPop_out(load_validBitDelay_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1__pushPop_out), .reset(load_reset));
  ShiftRegister_0_CEtrue_TY1 #(.INSTANCE_NAME("store_validBitDelay_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1_")) store_validBitDelay_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1_(.CLK(CLK), .CE(unnamedbinop12115USEDMULTIPLEbinop), .sr_input((1'd1)), .pushPop_out(store_validBitDelay_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1__pushPop_out));
endmodule

module incif_wrap648_inc8(input CLK, input CE, input [16:0] process_input, output [15:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] unnamedcast45USEDMULTIPLEcast = (process_input[15:0]);
  assign process_output = (((process_input[16]))?((({(unnamedcast45USEDMULTIPLEcast==(16'd648))})?((16'd0)):({(unnamedcast45USEDMULTIPLEcast+(16'd8))}))):(unnamedcast45USEDMULTIPLEcast));
  // function: process pure=true delay=0
endmodule

module RegBy_incif_wrap648_inc8_CEtrue_init0(input CLK, input set_valid, input CE, input [15:0] set_inp, input setby_valid, input setby_inp, output [15:0] SETBY_OUTPUT, output [15:0] GET_OUTPUT);
parameter INSTANCE_NAME="INST";
  reg [15:0] R = 16'd0;
  wire [15:0] regby_inner_process_output;
  always @(posedge CLK) begin if(set_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(setby_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,set_valid})+({4'b0,setby_valid})) > 5'd1) begin $display("error, function 'set' on instance 'R' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [16:0] unnamedcallArbitrate96USEDMULTIPLEcallArbitrate = {(set_valid||setby_valid),((set_valid)?(set_inp):(regby_inner_process_output))};
    always @ (posedge CLK) begin if ((unnamedcallArbitrate96USEDMULTIPLEcallArbitrate[16]) && CE) begin R <= (unnamedcallArbitrate96USEDMULTIPLEcallArbitrate[15:0]); end end
  assign SETBY_OUTPUT = regby_inner_process_output;
  assign GET_OUTPUT = R;
  // function: set pure=false ONLY WIRE
  // function: setby pure=false ONLY WIRE
  // function: get pure=true ONLY WIRE
  incif_wrap648_inc8 #(.INSTANCE_NAME("regby_inner")) regby_inner(.CLK(CLK), .CE(CE), .process_input({setby_inp,R}), .process_output(regby_inner_process_output));
endmodule

module incif_wrap482_incnil(input CLK, input CE, input [16:0] process_input, output [15:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] unnamedcast103USEDMULTIPLEcast = (process_input[15:0]);
  assign process_output = (((process_input[16]))?((({(unnamedcast103USEDMULTIPLEcast==(16'd482))})?((16'd0)):({(unnamedcast103USEDMULTIPLEcast+(16'd1))}))):(unnamedcast103USEDMULTIPLEcast));
  // function: process pure=true delay=0
endmodule

module RegBy_incif_wrap482_incnil_CEtrue_init0(input CLK, input set_valid, input CE, input [15:0] set_inp, input setby_valid, input setby_inp, output [15:0] SETBY_OUTPUT, output [15:0] GET_OUTPUT);
parameter INSTANCE_NAME="INST";
  reg [15:0] R = 16'd0;
  wire [15:0] regby_inner_process_output;
  always @(posedge CLK) begin if(set_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(setby_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,set_valid})+({4'b0,setby_valid})) > 5'd1) begin $display("error, function 'set' on instance 'R' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [16:0] unnamedcallArbitrate154USEDMULTIPLEcallArbitrate = {(set_valid||setby_valid),((set_valid)?(set_inp):(regby_inner_process_output))};
    always @ (posedge CLK) begin if ((unnamedcallArbitrate154USEDMULTIPLEcallArbitrate[16]) && CE) begin R <= (unnamedcallArbitrate154USEDMULTIPLEcallArbitrate[15:0]); end end
  assign SETBY_OUTPUT = regby_inner_process_output;
  assign GET_OUTPUT = R;
  // function: set pure=false ONLY WIRE
  // function: setby pure=false ONLY WIRE
  // function: get pure=true ONLY WIRE
  incif_wrap482_incnil #(.INSTANCE_NAME("regby_inner")) regby_inner(.CLK(CLK), .CE(CE), .process_input({setby_inp,R}), .process_output(regby_inner_process_output));
endmodule

module PadSeq_W640_H480_L8_R8_B1_Top1_T88(input CLK, output ready, input reset, input CE, input process_valid, input [63:0] process_input, output [64:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  wire [15:0] posX_padSeq_GET_OUTPUT;
  wire [15:0] unnamedcast166USEDMULTIPLEcast = (16'd648);
  wire [15:0] posY_padSeq_GET_OUTPUT;
  wire unnamedbinop178USEDMULTIPLEbinop = {({({((posX_padSeq_GET_OUTPUT)>=((16'd8)))}&&{((posX_padSeq_GET_OUTPUT)<(unnamedcast166USEDMULTIPLEcast))})}&&{({((posY_padSeq_GET_OUTPUT)>=((16'd1)))}&&{((posY_padSeq_GET_OUTPUT)<((16'd481)))})})};
  assign ready = unnamedbinop178USEDMULTIPLEbinop;
  reg [63:0] unnamedselect190_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect190_delay1_validunnamednull0_CECE <= ((unnamedbinop178USEDMULTIPLEbinop)?(process_input):({(8'd0),(8'd0),(8'd0),(8'd0),(8'd0),(8'd0),(8'd0),(8'd0)})); end end
  wire [15:0] posY_padSeq_SETBY_OUTPUT;
  wire [15:0] posX_padSeq_SETBY_OUTPUT;
  assign process_output = {(1'd1),unnamedselect190_delay1_validunnamednull0_CECE};
  // function: ready pure=true delay=0
  // function: reset pure=false delay=0
  // function: process pure=false delay=1
  RegBy_incif_wrap648_inc8_CEtrue_init0 #(.INSTANCE_NAME("posX_padSeq")) posX_padSeq(.CLK(CLK), .set_valid(reset), .CE(CE), .set_inp((16'd0)), .setby_valid(process_valid), .setby_inp((1'd1)), .SETBY_OUTPUT(posX_padSeq_SETBY_OUTPUT), .GET_OUTPUT(posX_padSeq_GET_OUTPUT));
  RegBy_incif_wrap482_incnil_CEtrue_init0 #(.INSTANCE_NAME("posY_padSeq")) posY_padSeq(.CLK(CLK), .set_valid(reset), .CE(CE), .set_inp((16'd0)), .setby_valid(process_valid), .setby_inp({(posX_padSeq_GET_OUTPUT==unnamedcast166USEDMULTIPLEcast)}), .SETBY_OUTPUT(posY_padSeq_SETBY_OUTPUT), .GET_OUTPUT(posY_padSeq_GET_OUTPUT));
endmodule

module WaitOnInput_PadSeq_W640_H480_L8_R8_B1_Top1_T88(input CLK, output ready, input reset, input CE, input process_valid, input [64:0] process_input, output [64:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  wire WaitOnInput_inner_ready;
  assign ready = WaitOnInput_inner_ready;
  wire unnamedbinop298USEDMULTIPLEbinop = {({({(~WaitOnInput_inner_ready)}||(process_input[64]))}&&process_valid)};
  wire [64:0] WaitOnInput_inner_process_output;
  reg unnamedbinop298_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedbinop298_delay1_validunnamednull0_CECE <= unnamedbinop298USEDMULTIPLEbinop; end end
  assign process_output = {{((WaitOnInput_inner_process_output[64])&&unnamedbinop298_delay1_validunnamednull0_CECE)},(WaitOnInput_inner_process_output[63:0])};
  // function: ready pure=true delay=0
  // function: reset pure=false delay=0
  // function: process pure=false delay=1
  PadSeq_W640_H480_L8_R8_B1_Top1_T88 #(.INSTANCE_NAME("WaitOnInput_inner")) WaitOnInput_inner(.CLK(CLK), .ready(WaitOnInput_inner_ready), .reset(reset), .CE(CE), .process_valid(unnamedbinop298USEDMULTIPLEbinop), .process_input((process_input[63:0])), .process_output(WaitOnInput_inner_process_output));
endmodule

module LiftHandshake_WaitOnInput_PadSeq_W640_H480_L8_R8_B1_Top1_T88(input CLK, input ready_downstream, output ready, input reset, input [64:0] process_input, output [64:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire inner_WaitOnInput_PadSeq_W640_H480_L8_R8_B1_Top1_T88_ready;
  assign ready = {(inner_WaitOnInput_PadSeq_W640_H480_L8_R8_B1_Top1_T88_ready&&ready_downstream)};
  wire unnamedbinop333USEDMULTIPLEbinop = {(reset||ready_downstream)};
  wire unnamedunary334USEDMULTIPLEunary = {(~reset)};
  wire [64:0] inner_WaitOnInput_PadSeq_W640_H480_L8_R8_B1_Top1_T88_process_output;
  wire validBitDelay_WaitOnInput_PadSeq_W640_H480_L8_R8_B1_Top1_T88_pushPop_out;
  wire [64:0] unnamedtuple366USEDMULTIPLEtuple = {{((inner_WaitOnInput_PadSeq_W640_H480_L8_R8_B1_Top1_T88_process_output[64])&&validBitDelay_WaitOnInput_PadSeq_W640_H480_L8_R8_B1_Top1_T88_pushPop_out)},(inner_WaitOnInput_PadSeq_W640_H480_L8_R8_B1_Top1_T88_process_output[63:0])};
  always @(posedge CLK) begin if({(~{((unnamedtuple366USEDMULTIPLEtuple[64])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: output valid bit should not be X!",INSTANCE_NAME); end end
  always @(posedge CLK) begin if({(~{((process_input[64])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = unnamedtuple366USEDMULTIPLEtuple;
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  WaitOnInput_PadSeq_W640_H480_L8_R8_B1_Top1_T88 #(.INSTANCE_NAME("inner_WaitOnInput_PadSeq_W640_H480_L8_R8_B1_Top1_T88")) inner_WaitOnInput_PadSeq_W640_H480_L8_R8_B1_Top1_T88(.CLK(CLK), .ready(inner_WaitOnInput_PadSeq_W640_H480_L8_R8_B1_Top1_T88_ready), .reset(reset), .CE(unnamedbinop333USEDMULTIPLEbinop), .process_valid(unnamedunary334USEDMULTIPLEunary), .process_input(process_input), .process_output(inner_WaitOnInput_PadSeq_W640_H480_L8_R8_B1_Top1_T88_process_output));
  ShiftRegister_1_CEtrue_TY1 #(.INSTANCE_NAME("validBitDelay_WaitOnInput_PadSeq_W640_H480_L8_R8_B1_Top1_T88")) validBitDelay_WaitOnInput_PadSeq_W640_H480_L8_R8_B1_Top1_T88(.CLK(CLK), .pushPop_valid(unnamedunary334USEDMULTIPLEunary), .CE(unnamedbinop333USEDMULTIPLEbinop), .sr_input((1'd1)), .pushPop_out(validBitDelay_WaitOnInput_PadSeq_W640_H480_L8_R8_B1_Top1_T88_pushPop_out), .reset(reset));
endmodule

module ShiftRegister_31_CEtrue_TY1(input CLK, input pushPop_valid, input CE, input sr_input, output pushPop_out, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'pushPop'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  reg SR31;
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR1' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR1' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR1' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6016USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(sr_input):((1'd0)))};
  reg SR1;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6016USEDMULTIPLEcallArbitrate[1]) && CE) begin SR1 <= (unnamedcallArbitrate6016USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR2' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR2' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR2' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6022USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR1):((1'd0)))};
  reg SR2;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6022USEDMULTIPLEcallArbitrate[1]) && CE) begin SR2 <= (unnamedcallArbitrate6022USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR3' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR3' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR3' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6028USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR2):((1'd0)))};
  reg SR3;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6028USEDMULTIPLEcallArbitrate[1]) && CE) begin SR3 <= (unnamedcallArbitrate6028USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR4' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR4' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR4' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6034USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR3):((1'd0)))};
  reg SR4;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6034USEDMULTIPLEcallArbitrate[1]) && CE) begin SR4 <= (unnamedcallArbitrate6034USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR5' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR5' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR5' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6040USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR4):((1'd0)))};
  reg SR5;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6040USEDMULTIPLEcallArbitrate[1]) && CE) begin SR5 <= (unnamedcallArbitrate6040USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR6' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR6' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR6' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6046USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR5):((1'd0)))};
  reg SR6;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6046USEDMULTIPLEcallArbitrate[1]) && CE) begin SR6 <= (unnamedcallArbitrate6046USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR7' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR7' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR7' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6052USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR6):((1'd0)))};
  reg SR7;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6052USEDMULTIPLEcallArbitrate[1]) && CE) begin SR7 <= (unnamedcallArbitrate6052USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR8' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR8' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR8' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6058USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR7):((1'd0)))};
  reg SR8;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6058USEDMULTIPLEcallArbitrate[1]) && CE) begin SR8 <= (unnamedcallArbitrate6058USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR9' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR9' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR9' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6064USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR8):((1'd0)))};
  reg SR9;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6064USEDMULTIPLEcallArbitrate[1]) && CE) begin SR9 <= (unnamedcallArbitrate6064USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR10' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR10' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR10' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6070USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR9):((1'd0)))};
  reg SR10;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6070USEDMULTIPLEcallArbitrate[1]) && CE) begin SR10 <= (unnamedcallArbitrate6070USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR11' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR11' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR11' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6076USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR10):((1'd0)))};
  reg SR11;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6076USEDMULTIPLEcallArbitrate[1]) && CE) begin SR11 <= (unnamedcallArbitrate6076USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR12' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR12' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR12' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6082USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR11):((1'd0)))};
  reg SR12;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6082USEDMULTIPLEcallArbitrate[1]) && CE) begin SR12 <= (unnamedcallArbitrate6082USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR13' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR13' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR13' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6088USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR12):((1'd0)))};
  reg SR13;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6088USEDMULTIPLEcallArbitrate[1]) && CE) begin SR13 <= (unnamedcallArbitrate6088USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR14' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR14' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR14' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6094USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR13):((1'd0)))};
  reg SR14;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6094USEDMULTIPLEcallArbitrate[1]) && CE) begin SR14 <= (unnamedcallArbitrate6094USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR15' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR15' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR15' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6100USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR14):((1'd0)))};
  reg SR15;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6100USEDMULTIPLEcallArbitrate[1]) && CE) begin SR15 <= (unnamedcallArbitrate6100USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR16' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR16' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR16' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6106USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR15):((1'd0)))};
  reg SR16;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6106USEDMULTIPLEcallArbitrate[1]) && CE) begin SR16 <= (unnamedcallArbitrate6106USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR17' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR17' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR17' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6112USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR16):((1'd0)))};
  reg SR17;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6112USEDMULTIPLEcallArbitrate[1]) && CE) begin SR17 <= (unnamedcallArbitrate6112USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR18' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR18' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR18' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6118USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR17):((1'd0)))};
  reg SR18;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6118USEDMULTIPLEcallArbitrate[1]) && CE) begin SR18 <= (unnamedcallArbitrate6118USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR19' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR19' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR19' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6124USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR18):((1'd0)))};
  reg SR19;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6124USEDMULTIPLEcallArbitrate[1]) && CE) begin SR19 <= (unnamedcallArbitrate6124USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR20' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR20' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR20' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6130USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR19):((1'd0)))};
  reg SR20;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6130USEDMULTIPLEcallArbitrate[1]) && CE) begin SR20 <= (unnamedcallArbitrate6130USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR21' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR21' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR21' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6136USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR20):((1'd0)))};
  reg SR21;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6136USEDMULTIPLEcallArbitrate[1]) && CE) begin SR21 <= (unnamedcallArbitrate6136USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR22' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR22' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR22' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6142USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR21):((1'd0)))};
  reg SR22;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6142USEDMULTIPLEcallArbitrate[1]) && CE) begin SR22 <= (unnamedcallArbitrate6142USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR23' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR23' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR23' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6148USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR22):((1'd0)))};
  reg SR23;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6148USEDMULTIPLEcallArbitrate[1]) && CE) begin SR23 <= (unnamedcallArbitrate6148USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR24' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR24' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR24' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6154USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR23):((1'd0)))};
  reg SR24;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6154USEDMULTIPLEcallArbitrate[1]) && CE) begin SR24 <= (unnamedcallArbitrate6154USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR25' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR25' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR25' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6160USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR24):((1'd0)))};
  reg SR25;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6160USEDMULTIPLEcallArbitrate[1]) && CE) begin SR25 <= (unnamedcallArbitrate6160USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR26' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR26' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR26' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6166USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR25):((1'd0)))};
  reg SR26;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6166USEDMULTIPLEcallArbitrate[1]) && CE) begin SR26 <= (unnamedcallArbitrate6166USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR27' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR27' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR27' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6172USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR26):((1'd0)))};
  reg SR27;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6172USEDMULTIPLEcallArbitrate[1]) && CE) begin SR27 <= (unnamedcallArbitrate6172USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR28' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR28' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR28' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6178USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR27):((1'd0)))};
  reg SR28;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6178USEDMULTIPLEcallArbitrate[1]) && CE) begin SR28 <= (unnamedcallArbitrate6178USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR29' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR29' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR29' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6184USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR28):((1'd0)))};
  reg SR29;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6184USEDMULTIPLEcallArbitrate[1]) && CE) begin SR29 <= (unnamedcallArbitrate6184USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR30' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR30' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR30' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6190USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR29):((1'd0)))};
  reg SR30;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6190USEDMULTIPLEcallArbitrate[1]) && CE) begin SR30 <= (unnamedcallArbitrate6190USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR31' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR31' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR31' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6196USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR30):((1'd0)))};
    always @ (posedge CLK) begin if ((unnamedcallArbitrate6196USEDMULTIPLEcallArbitrate[1]) && CE) begin SR31 <= (unnamedcallArbitrate6196USEDMULTIPLEcallArbitrate[0]); end end
  assign pushPop_out = SR31;
  // function: pushPop pure=false delay=0
  // function: reset pure=false delay=0
endmodule

module blackLevel(input CLK, input process_CE, input [7:0] blInput, output [7:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [8:0] unnamedcast2066 = {1'b0,blInput}; // wire for int size extend (cast)
  wire [8:0] unnamedcast2068 = {1'b0,(8'd90)}; // wire for int size extend (cast)
  wire [9:0] unnamedcast2069 = { {1{unnamedcast2066[8]}},unnamedcast2066[8:0]};// wire for $signed
  wire [9:0] unnamedcast2070 = { {1{unnamedcast2068[8]}},unnamedcast2068[8:0]};// wire for $signed
  reg [9:0] unnamedbinop2071_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2071_delay1_validunnamednull0_CEprocess_CE <= {($signed(unnamedcast2069)-$signed(unnamedcast2070))}; end end
  wire [8:0] unnamedcast2073 = {1'b0,(8'd197)}; // wire for int size extend (cast)
  reg [18:0] unnamedcast2075_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2075_delay1_validunnamednull0_CEprocess_CE <= { {10{unnamedcast2073[8]}},unnamedcast2073[8:0]}; end end
  wire [18:0] unnamedcast2074 = { {9{unnamedbinop2071_delay1_validunnamednull0_CEprocess_CE[9]}},unnamedbinop2071_delay1_validunnamednull0_CEprocess_CE[9:0]};// wire for $signed
  reg [18:0] unnamedbinop2076_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2076_delay1_validunnamednull0_CEprocess_CE <= {($signed(unnamedcast2074)*$signed(unnamedcast2075_delay1_validunnamednull0_CEprocess_CE))}; end end
  reg [18:0] unnamedunary2077_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedunary2077_delay1_validunnamednull0_CEprocess_CE <= {((unnamedbinop2076_delay1_validunnamednull0_CEprocess_CE[18])?(-unnamedbinop2076_delay1_validunnamednull0_CEprocess_CE):(unnamedbinop2076_delay1_validunnamednull0_CEprocess_CE))}; end end
  reg [18:0] unnamedcast2080_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2080_delay1_validunnamednull0_CEprocess_CE <= (19'd7); end end
  reg [18:0] unnamedcast2080_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2080_delay2_validunnamednull0_CEprocess_CE <= unnamedcast2080_delay1_validunnamednull0_CEprocess_CE; end end
  reg [18:0] unnamedcast2080_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2080_delay3_validunnamednull0_CEprocess_CE <= unnamedcast2080_delay2_validunnamednull0_CEprocess_CE; end end
  reg [18:0] unnamedbinop2081_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2081_delay1_validunnamednull0_CEprocess_CE <= {(unnamedunary2077_delay1_validunnamednull0_CEprocess_CE>>>unnamedcast2080_delay3_validunnamednull0_CEprocess_CE)}; end end
  wire [11:0] unnamedcast2082USEDMULTIPLEcast = unnamedbinop2081_delay1_validunnamednull0_CEprocess_CE[11:0];
  reg [11:0] unnamedcast2084_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2084_delay1_validunnamednull0_CEprocess_CE <= {4'b0,(8'd255)}; end end
  reg [11:0] unnamedcast2084_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2084_delay2_validunnamednull0_CEprocess_CE <= unnamedcast2084_delay1_validunnamednull0_CEprocess_CE; end end
  reg [11:0] unnamedcast2084_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2084_delay3_validunnamednull0_CEprocess_CE <= unnamedcast2084_delay2_validunnamednull0_CEprocess_CE; end end
  reg [11:0] unnamedcast2084_delay4_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2084_delay4_validunnamednull0_CEprocess_CE <= unnamedcast2084_delay3_validunnamednull0_CEprocess_CE; end end
  reg unnamedbinop2085_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2085_delay1_validunnamednull0_CEprocess_CE <= {((unnamedcast2082USEDMULTIPLEcast)>(unnamedcast2084_delay4_validunnamednull0_CEprocess_CE))}; end end
  reg [11:0] unnamedcast2087_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2087_delay1_validunnamednull0_CEprocess_CE <= (12'd255); end end
  reg [11:0] unnamedcast2087_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2087_delay2_validunnamednull0_CEprocess_CE <= unnamedcast2087_delay1_validunnamednull0_CEprocess_CE; end end
  reg [11:0] unnamedcast2087_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2087_delay3_validunnamednull0_CEprocess_CE <= unnamedcast2087_delay2_validunnamednull0_CEprocess_CE; end end
  reg [11:0] unnamedcast2087_delay4_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2087_delay4_validunnamednull0_CEprocess_CE <= unnamedcast2087_delay3_validunnamednull0_CEprocess_CE; end end
  reg [11:0] unnamedcast2087_delay5_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2087_delay5_validunnamednull0_CEprocess_CE <= unnamedcast2087_delay4_validunnamednull0_CEprocess_CE; end end
  reg [11:0] unnamedcast2082_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2082_delay1_validunnamednull0_CEprocess_CE <= unnamedcast2082USEDMULTIPLEcast; end end
  reg [11:0] unnamedselect2088_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedselect2088_delay1_validunnamednull0_CEprocess_CE <= ((unnamedbinop2085_delay1_validunnamednull0_CEprocess_CE)?(unnamedcast2087_delay5_validunnamednull0_CEprocess_CE):(unnamedcast2082_delay1_validunnamednull0_CEprocess_CE)); end end
  assign process_output = unnamedselect2088_delay1_validunnamednull0_CEprocess_CE[7:0];
  // function: process pure=true delay=6
endmodule

module map_blackLevel_W8_H1(input CLK, input process_CE, input [63:0] process_input, output [63:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [7:0] inner0_0_process_output;
  wire [7:0] inner1_0_process_output;
  wire [7:0] inner2_0_process_output;
  wire [7:0] inner3_0_process_output;
  wire [7:0] inner4_0_process_output;
  wire [7:0] inner5_0_process_output;
  wire [7:0] inner6_0_process_output;
  wire [7:0] inner7_0_process_output;
  assign process_output = {inner7_0_process_output,inner6_0_process_output,inner5_0_process_output,inner4_0_process_output,inner3_0_process_output,inner2_0_process_output,inner1_0_process_output,inner0_0_process_output};
  // function: process pure=true delay=6
  blackLevel #(.INSTANCE_NAME("inner0_0")) inner0_0(.CLK(CLK), .process_CE(process_CE), .blInput(({process_input[7:0]})), .process_output(inner0_0_process_output));
  blackLevel #(.INSTANCE_NAME("inner1_0")) inner1_0(.CLK(CLK), .process_CE(process_CE), .blInput(({process_input[15:8]})), .process_output(inner1_0_process_output));
  blackLevel #(.INSTANCE_NAME("inner2_0")) inner2_0(.CLK(CLK), .process_CE(process_CE), .blInput(({process_input[23:16]})), .process_output(inner2_0_process_output));
  blackLevel #(.INSTANCE_NAME("inner3_0")) inner3_0(.CLK(CLK), .process_CE(process_CE), .blInput(({process_input[31:24]})), .process_output(inner3_0_process_output));
  blackLevel #(.INSTANCE_NAME("inner4_0")) inner4_0(.CLK(CLK), .process_CE(process_CE), .blInput(({process_input[39:32]})), .process_output(inner4_0_process_output));
  blackLevel #(.INSTANCE_NAME("inner5_0")) inner5_0(.CLK(CLK), .process_CE(process_CE), .blInput(({process_input[47:40]})), .process_output(inner5_0_process_output));
  blackLevel #(.INSTANCE_NAME("inner6_0")) inner6_0(.CLK(CLK), .process_CE(process_CE), .blInput(({process_input[55:48]})), .process_output(inner6_0_process_output));
  blackLevel #(.INSTANCE_NAME("inner7_0")) inner7_0(.CLK(CLK), .process_CE(process_CE), .blInput(({process_input[63:56]})), .process_output(inner7_0_process_output));
endmodule

module incif_wrap81_incnil(input CLK, input CE, input [16:0] process_input, output [15:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] unnamedcast4082USEDMULTIPLEcast = (process_input[15:0]);
  assign process_output = (((process_input[16]))?((({(unnamedcast4082USEDMULTIPLEcast==(16'd81))})?((16'd0)):({(unnamedcast4082USEDMULTIPLEcast+(16'd1))}))):(unnamedcast4082USEDMULTIPLEcast));
  // function: process pure=true delay=0
endmodule

module RegBy_incif_wrap81_incnil_CEtrue_initnil(input CLK, input set_valid, input CE, input [15:0] set_inp, input setby_valid, input setby_inp, output [15:0] SETBY_OUTPUT, output [15:0] GET_OUTPUT);
parameter INSTANCE_NAME="INST";
  reg [15:0] R;
  wire [15:0] regby_inner_process_output;
  always @(posedge CLK) begin if(set_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(setby_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,set_valid})+({4'b0,setby_valid})) > 5'd1) begin $display("error, function 'set' on instance 'R' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [16:0] unnamedcallArbitrate4133USEDMULTIPLEcallArbitrate = {(set_valid||setby_valid),((set_valid)?(set_inp):(regby_inner_process_output))};
    always @ (posedge CLK) begin if ((unnamedcallArbitrate4133USEDMULTIPLEcallArbitrate[16]) && CE) begin R <= (unnamedcallArbitrate4133USEDMULTIPLEcallArbitrate[15:0]); end end
  assign SETBY_OUTPUT = regby_inner_process_output;
  assign GET_OUTPUT = R;
  // function: set pure=false ONLY WIRE
  // function: setby pure=false ONLY WIRE
  // function: get pure=true ONLY WIRE
  incif_wrap81_incnil #(.INSTANCE_NAME("regby_inner")) regby_inner(.CLK(CLK), .CE(CE), .process_input({setby_inp,R}), .process_output(regby_inner_process_output));
endmodule

module bramSDP_WAROtrue_size1024_bw8_obwnil_CEtrue_inittable__0x422b92d8(input CLK, input writeAndReturnOriginal_valid, input writeAndReturnOriginal_CE, input [70:0] inp, output [63:0] WARO_OUT);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(writeAndReturnOriginal_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'writeAndReturnOriginal'", INSTANCE_NAME);  end end
  wire [8:0] unnamedcast4144USEDMULTIPLEcast = {2'b0,(inp[6:0])};
  wire [63:0] unnamedcast4142USEDMULTIPLEcast = (inp[70:7]);
  wire [31:0] bram_0_SET_AND_RETURN_ORIG_OUTPUT;
  wire [31:0] bram_1_SET_AND_RETURN_ORIG_OUTPUT;
  assign WARO_OUT = {bram_1_SET_AND_RETURN_ORIG_OUTPUT,bram_0_SET_AND_RETURN_ORIG_OUTPUT};
  // function: writeAndReturnOriginal pure=false delay=1
  reg [31:0] bram_0_DI_B;
reg [8:0] bram_0_addr_B;
wire [31:0] bram_0_DO_B;
wire [40:0] bram_0_INPUT;
assign bram_0_INPUT = {unnamedcast4142USEDMULTIPLEcast[31:0],unnamedcast4144USEDMULTIPLEcast};
RAMB16_S36_S36 #(.WRITE_MODE_A("READ_FIRST"),.WRITE_MODE_B("READ_FIRST"),.INIT_00(256'h1f1e1d1c1b1a191817161514131211100f0e0d0c0b0a09080706050403020100),.INIT_01(256'h3f3e3d3c3b3a393837363534333231302f2e2d2c2b2a29282726252423222120),.INIT_02(256'h5f5e5d5c5b5a595857565554535251504f4e4d4c4b4a49484746454443424140),.INIT_03(256'h7f7e7d7c7b7a797877767574737271706f6e6d6c6b6a69686766656463626160),.INIT_04(256'h9f9e9d9c9b9a999897969594939291908f8e8d8c8b8a89888786858483828180),.INIT_05(256'hbfbebdbcbbbab9b8b7b6b5b4b3b2b1b0afaeadacabaaa9a8a7a6a5a4a3a2a1a0),.INIT_06(256'hdfdedddcdbdad9d8d7d6d5d4d3d2d1d0cfcecdcccbcac9c8c7c6c5c4c3c2c1c0),.INIT_07(256'hfffefdfcfbfaf9f8f7f6f5f4f3f2f1f0efeeedecebeae9e8e7e6e5e4e3e2e1e0),.INIT_08(256'h1f1e1d1c1b1a191817161514131211100f0e0d0c0b0a09080706050403020100),.INIT_09(256'h3f3e3d3c3b3a393837363534333231302f2e2d2c2b2a29282726252423222120),.INIT_0A(256'h5f5e5d5c5b5a595857565554535251504f4e4d4c4b4a49484746454443424140),.INIT_0B(256'h7f7e7d7c7b7a797877767574737271706f6e6d6c6b6a69686766656463626160),.INIT_0C(256'h9f9e9d9c9b9a999897969594939291908f8e8d8c8b8a89888786858483828180),.INIT_0D(256'hbfbebdbcbbbab9b8b7b6b5b4b3b2b1b0afaeadacabaaa9a8a7a6a5a4a3a2a1a0),.INIT_0E(256'hdfdedddcdbdad9d8d7d6d5d4d3d2d1d0cfcecdcccbcac9c8c7c6c5c4c3c2c1c0),.INIT_0F(256'hfffefdfcfbfaf9f8f7f6f5f4f3f2f1f0efeeedecebeae9e8e7e6e5e4e3e2e1e0),.INIT_10(256'h1f1e1d1c1b1a191817161514131211100f0e0d0c0b0a09080706050403020100),.INIT_11(256'h3f3e3d3c3b3a393837363534333231302f2e2d2c2b2a29282726252423222120),.INIT_12(256'h5f5e5d5c5b5a595857565554535251504f4e4d4c4b4a49484746454443424140),.INIT_13(256'h7f7e7d7c7b7a797877767574737271706f6e6d6c6b6a69686766656463626160),.INIT_14(256'h9f9e9d9c9b9a999897969594939291908f8e8d8c8b8a89888786858483828180),.INIT_15(256'hbfbebdbcbbbab9b8b7b6b5b4b3b2b1b0afaeadacabaaa9a8a7a6a5a4a3a2a1a0),.INIT_16(256'hdfdedddcdbdad9d8d7d6d5d4d3d2d1d0cfcecdcccbcac9c8c7c6c5c4c3c2c1c0),.INIT_17(256'hfffefdfcfbfaf9f8f7f6f5f4f3f2f1f0efeeedecebeae9e8e7e6e5e4e3e2e1e0),.INIT_18(256'h1f1e1d1c1b1a191817161514131211100f0e0d0c0b0a09080706050403020100),.INIT_19(256'h3f3e3d3c3b3a393837363534333231302f2e2d2c2b2a29282726252423222120),.INIT_1A(256'h5f5e5d5c5b5a595857565554535251504f4e4d4c4b4a49484746454443424140),.INIT_1B(256'h7f7e7d7c7b7a797877767574737271706f6e6d6c6b6a69686766656463626160),.INIT_1C(256'h9f9e9d9c9b9a999897969594939291908f8e8d8c8b8a89888786858483828180),.INIT_1D(256'hbfbebdbcbbbab9b8b7b6b5b4b3b2b1b0afaeadacabaaa9a8a7a6a5a4a3a2a1a0),.INIT_1E(256'hdfdedddcdbdad9d8d7d6d5d4d3d2d1d0cfcecdcccbcac9c8c7c6c5c4c3c2c1c0),.INIT_1F(256'hfffefdfcfbfaf9f8f7f6f5f4f3f2f1f0efeeedecebeae9e8e7e6e5e4e3e2e1e0),.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)) bram_0 (
.DIPA(4'b0),
.DIPB(4'b0),
.DIA(bram_0_INPUT[40:9]),
.DIB(bram_0_DI_B),
.DOA(bram_0_SET_AND_RETURN_ORIG_OUTPUT),
.DOB(bram_0_DO_B),
.ADDRA(bram_0_INPUT[8:0]),
.ADDRB(bram_0_addr_B),
.WEA(writeAndReturnOriginal_valid),
.WEB(1'd0),
.ENA(writeAndReturnOriginal_CE),
.ENB(writeAndReturnOriginal_CE),
.CLKA(CLK),
.CLKB(CLK),
.SSRA(1'b0),
.SSRB(1'b0)
);


  reg [31:0] bram_1_DI_B;
reg [8:0] bram_1_addr_B;
wire [31:0] bram_1_DO_B;
wire [40:0] bram_1_INPUT;
assign bram_1_INPUT = {unnamedcast4142USEDMULTIPLEcast[63:32],unnamedcast4144USEDMULTIPLEcast};
RAMB16_S36_S36 #(.WRITE_MODE_A("READ_FIRST"),.WRITE_MODE_B("READ_FIRST"),.INIT_00(256'h1f1e1d1c1b1a191817161514131211100f0e0d0c0b0a09080706050403020100),.INIT_01(256'h3f3e3d3c3b3a393837363534333231302f2e2d2c2b2a29282726252423222120),.INIT_02(256'h5f5e5d5c5b5a595857565554535251504f4e4d4c4b4a49484746454443424140),.INIT_03(256'h7f7e7d7c7b7a797877767574737271706f6e6d6c6b6a69686766656463626160),.INIT_04(256'h9f9e9d9c9b9a999897969594939291908f8e8d8c8b8a89888786858483828180),.INIT_05(256'hbfbebdbcbbbab9b8b7b6b5b4b3b2b1b0afaeadacabaaa9a8a7a6a5a4a3a2a1a0),.INIT_06(256'hdfdedddcdbdad9d8d7d6d5d4d3d2d1d0cfcecdcccbcac9c8c7c6c5c4c3c2c1c0),.INIT_07(256'hfffefdfcfbfaf9f8f7f6f5f4f3f2f1f0efeeedecebeae9e8e7e6e5e4e3e2e1e0),.INIT_08(256'h1f1e1d1c1b1a191817161514131211100f0e0d0c0b0a09080706050403020100),.INIT_09(256'h3f3e3d3c3b3a393837363534333231302f2e2d2c2b2a29282726252423222120),.INIT_0A(256'h5f5e5d5c5b5a595857565554535251504f4e4d4c4b4a49484746454443424140),.INIT_0B(256'h7f7e7d7c7b7a797877767574737271706f6e6d6c6b6a69686766656463626160),.INIT_0C(256'h9f9e9d9c9b9a999897969594939291908f8e8d8c8b8a89888786858483828180),.INIT_0D(256'hbfbebdbcbbbab9b8b7b6b5b4b3b2b1b0afaeadacabaaa9a8a7a6a5a4a3a2a1a0),.INIT_0E(256'hdfdedddcdbdad9d8d7d6d5d4d3d2d1d0cfcecdcccbcac9c8c7c6c5c4c3c2c1c0),.INIT_0F(256'hfffefdfcfbfaf9f8f7f6f5f4f3f2f1f0efeeedecebeae9e8e7e6e5e4e3e2e1e0),.INIT_10(256'h1f1e1d1c1b1a191817161514131211100f0e0d0c0b0a09080706050403020100),.INIT_11(256'h3f3e3d3c3b3a393837363534333231302f2e2d2c2b2a29282726252423222120),.INIT_12(256'h5f5e5d5c5b5a595857565554535251504f4e4d4c4b4a49484746454443424140),.INIT_13(256'h7f7e7d7c7b7a797877767574737271706f6e6d6c6b6a69686766656463626160),.INIT_14(256'h9f9e9d9c9b9a999897969594939291908f8e8d8c8b8a89888786858483828180),.INIT_15(256'hbfbebdbcbbbab9b8b7b6b5b4b3b2b1b0afaeadacabaaa9a8a7a6a5a4a3a2a1a0),.INIT_16(256'hdfdedddcdbdad9d8d7d6d5d4d3d2d1d0cfcecdcccbcac9c8c7c6c5c4c3c2c1c0),.INIT_17(256'hfffefdfcfbfaf9f8f7f6f5f4f3f2f1f0efeeedecebeae9e8e7e6e5e4e3e2e1e0),.INIT_18(256'h1f1e1d1c1b1a191817161514131211100f0e0d0c0b0a09080706050403020100),.INIT_19(256'h3f3e3d3c3b3a393837363534333231302f2e2d2c2b2a29282726252423222120),.INIT_1A(256'h5f5e5d5c5b5a595857565554535251504f4e4d4c4b4a49484746454443424140),.INIT_1B(256'h7f7e7d7c7b7a797877767574737271706f6e6d6c6b6a69686766656463626160),.INIT_1C(256'h9f9e9d9c9b9a999897969594939291908f8e8d8c8b8a89888786858483828180),.INIT_1D(256'hbfbebdbcbbbab9b8b7b6b5b4b3b2b1b0afaeadacabaaa9a8a7a6a5a4a3a2a1a0),.INIT_1E(256'hdfdedddcdbdad9d8d7d6d5d4d3d2d1d0cfcecdcccbcac9c8c7c6c5c4c3c2c1c0),.INIT_1F(256'hfffefdfcfbfaf9f8f7f6f5f4f3f2f1f0efeeedecebeae9e8e7e6e5e4e3e2e1e0),.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)) bram_1 (
.DIPA(4'b0),
.DIPB(4'b0),
.DIA(bram_1_INPUT[40:9]),
.DIB(bram_1_DI_B),
.DOA(bram_1_SET_AND_RETURN_ORIG_OUTPUT),
.DOB(bram_1_DO_B),
.ADDRA(bram_1_INPUT[8:0]),
.ADDRB(bram_1_addr_B),
.WEA(writeAndReturnOriginal_valid),
.WEB(1'd0),
.ENA(writeAndReturnOriginal_CE),
.ENB(writeAndReturnOriginal_CE),
.CLKA(CLK),
.CLKB(CLK),
.SSRA(1'b0),
.SSRB(1'b0)
);


endmodule

module linebuffer_w656_h482_T8_ymin_2_Auint8(input CLK, input process_valid, input CE, input [63:0] process_input, output [191:0] process_output, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  wire [15:0] addr_GET_OUTPUT;
  wire [6:0] unnamedcast4220USEDMULTIPLEcast = addr_GET_OUTPUT[6:0];
  reg [6:0] unnamedcast4220_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4220_delay1_validunnamednull0_CECE <= unnamedcast4220USEDMULTIPLEcast; end end
  wire [63:0] lb_m0_WARO_OUT;
  wire [63:0] unnamedcast4200USEDMULTIPLEcast = lb_m0_WARO_OUT[63:0];
  reg process_valid_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay1_validunnamednull0_CECE <= process_valid; end end
  wire [63:0] lb_m1_WARO_OUT;
  wire [63:0] unnamedcast4224USEDMULTIPLEcast = lb_m1_WARO_OUT[63:0];
  reg [7:0] unnamedcast4202_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4202_delay1_validunnamednull0_CECE <= ({unnamedcast4200USEDMULTIPLEcast[7:0]}); end end
  reg [7:0] unnamedcast4204_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4204_delay1_validunnamednull0_CECE <= ({unnamedcast4200USEDMULTIPLEcast[15:8]}); end end
  reg [7:0] unnamedcast4206_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4206_delay1_validunnamednull0_CECE <= ({unnamedcast4200USEDMULTIPLEcast[23:16]}); end end
  reg [7:0] unnamedcast4208_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4208_delay1_validunnamednull0_CECE <= ({unnamedcast4200USEDMULTIPLEcast[31:24]}); end end
  reg [7:0] unnamedcast4210_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4210_delay1_validunnamednull0_CECE <= ({unnamedcast4200USEDMULTIPLEcast[39:32]}); end end
  reg [7:0] unnamedcast4212_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4212_delay1_validunnamednull0_CECE <= ({unnamedcast4200USEDMULTIPLEcast[47:40]}); end end
  reg [7:0] unnamedcast4214_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4214_delay1_validunnamednull0_CECE <= ({unnamedcast4200USEDMULTIPLEcast[55:48]}); end end
  reg [7:0] unnamedcast4216_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4216_delay1_validunnamednull0_CECE <= ({unnamedcast4200USEDMULTIPLEcast[63:56]}); end end
  reg [7:0] unnamedcast4154_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4154_delay1_validunnamednull0_CECE <= ({process_input[7:0]}); end end
  reg [7:0] unnamedcast4154_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4154_delay2_validunnamednull0_CECE <= unnamedcast4154_delay1_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast4156_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4156_delay1_validunnamednull0_CECE <= ({process_input[15:8]}); end end
  reg [7:0] unnamedcast4156_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4156_delay2_validunnamednull0_CECE <= unnamedcast4156_delay1_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast4158_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4158_delay1_validunnamednull0_CECE <= ({process_input[23:16]}); end end
  reg [7:0] unnamedcast4158_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4158_delay2_validunnamednull0_CECE <= unnamedcast4158_delay1_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast4160_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4160_delay1_validunnamednull0_CECE <= ({process_input[31:24]}); end end
  reg [7:0] unnamedcast4160_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4160_delay2_validunnamednull0_CECE <= unnamedcast4160_delay1_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast4162_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4162_delay1_validunnamednull0_CECE <= ({process_input[39:32]}); end end
  reg [7:0] unnamedcast4162_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4162_delay2_validunnamednull0_CECE <= unnamedcast4162_delay1_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast4164_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4164_delay1_validunnamednull0_CECE <= ({process_input[47:40]}); end end
  reg [7:0] unnamedcast4164_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4164_delay2_validunnamednull0_CECE <= unnamedcast4164_delay1_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast4166_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4166_delay1_validunnamednull0_CECE <= ({process_input[55:48]}); end end
  reg [7:0] unnamedcast4166_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4166_delay2_validunnamednull0_CECE <= unnamedcast4166_delay1_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast4168_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4168_delay1_validunnamednull0_CECE <= ({process_input[63:56]}); end end
  reg [7:0] unnamedcast4168_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast4168_delay2_validunnamednull0_CECE <= unnamedcast4168_delay1_validunnamednull0_CECE; end end
  wire [15:0] addr_SETBY_OUTPUT;
  assign process_output = {unnamedcast4168_delay2_validunnamednull0_CECE,unnamedcast4166_delay2_validunnamednull0_CECE,unnamedcast4164_delay2_validunnamednull0_CECE,unnamedcast4162_delay2_validunnamednull0_CECE,unnamedcast4160_delay2_validunnamednull0_CECE,unnamedcast4158_delay2_validunnamednull0_CECE,unnamedcast4156_delay2_validunnamednull0_CECE,unnamedcast4154_delay2_validunnamednull0_CECE,unnamedcast4216_delay1_validunnamednull0_CECE,unnamedcast4214_delay1_validunnamednull0_CECE,unnamedcast4212_delay1_validunnamednull0_CECE,unnamedcast4210_delay1_validunnamednull0_CECE,unnamedcast4208_delay1_validunnamednull0_CECE,unnamedcast4206_delay1_validunnamednull0_CECE,unnamedcast4204_delay1_validunnamednull0_CECE,unnamedcast4202_delay1_validunnamednull0_CECE,({unnamedcast4224USEDMULTIPLEcast[63:56]}),({unnamedcast4224USEDMULTIPLEcast[55:48]}),({unnamedcast4224USEDMULTIPLEcast[47:40]}),({unnamedcast4224USEDMULTIPLEcast[39:32]}),({unnamedcast4224USEDMULTIPLEcast[31:24]}),({unnamedcast4224USEDMULTIPLEcast[23:16]}),({unnamedcast4224USEDMULTIPLEcast[15:8]}),({unnamedcast4224USEDMULTIPLEcast[7:0]})};
  // function: process pure=false delay=2
  // function: reset pure=false delay=0
  RegBy_incif_wrap81_incnil_CEtrue_initnil #(.INSTANCE_NAME("addr")) addr(.CLK(CLK), .set_valid(reset), .CE(CE), .set_inp((16'd0)), .setby_valid(process_valid), .setby_inp((1'd1)), .SETBY_OUTPUT(addr_SETBY_OUTPUT), .GET_OUTPUT(addr_GET_OUTPUT));
  bramSDP_WAROtrue_size1024_bw8_obwnil_CEtrue_inittable__0x422b92d8 #(.INSTANCE_NAME("lb_m0")) lb_m0(.CLK(CLK), .writeAndReturnOriginal_valid(process_valid), .writeAndReturnOriginal_CE(CE), .inp({process_input,unnamedcast4220USEDMULTIPLEcast}), .WARO_OUT(lb_m0_WARO_OUT));
  bramSDP_WAROtrue_size1024_bw8_obwnil_CEtrue_inittable__0x422b92d8 #(.INSTANCE_NAME("lb_m1")) lb_m1(.CLK(CLK), .writeAndReturnOriginal_valid(process_valid_delay1_validunnamednull0_CECE), .writeAndReturnOriginal_CE(CE), .inp({unnamedcast4200USEDMULTIPLEcast,unnamedcast4220_delay1_validunnamednull0_CECE}), .WARO_OUT(lb_m1_WARO_OUT));
endmodule

module SSR_W3_H3_T8_Auint8(input CLK, input process_valid, input process_CE, input [191:0] inp, output [239:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  reg [7:0] SR_x0_y0;
  reg [7:0] SR_x1_y0;
  wire [7:0] unnamedcast4010USEDMULTIPLEcast = ({inp[55:48]});
  wire [7:0] unnamedcast4008USEDMULTIPLEcast = ({inp[63:56]});
  reg [7:0] SR_x0_y1;
  reg [7:0] SR_x1_y1;
  wire [7:0] unnamedcast4034USEDMULTIPLEcast = ({inp[119:112]});
  wire [7:0] unnamedcast4032USEDMULTIPLEcast = ({inp[127:120]});
  reg [7:0] SR_x0_y2;
  reg [7:0] SR_x1_y2;
  wire [7:0] unnamedcast4058USEDMULTIPLEcast = ({inp[183:176]});
  wire [7:0] unnamedcast4056USEDMULTIPLEcast = ({inp[191:184]});
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x1_y0 <= unnamedcast4008USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x0_y0 <= unnamedcast4010USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x1_y1 <= unnamedcast4032USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x0_y1 <= unnamedcast4034USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x1_y2 <= unnamedcast4056USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x0_y2 <= unnamedcast4058USEDMULTIPLEcast; end end
  assign process_output = {unnamedcast4056USEDMULTIPLEcast,unnamedcast4058USEDMULTIPLEcast,({inp[175:168]}),({inp[167:160]}),({inp[159:152]}),({inp[151:144]}),({inp[143:136]}),({inp[135:128]}),SR_x1_y2,SR_x0_y2,unnamedcast4032USEDMULTIPLEcast,unnamedcast4034USEDMULTIPLEcast,({inp[111:104]}),({inp[103:96]}),({inp[95:88]}),({inp[87:80]}),({inp[79:72]}),({inp[71:64]}),SR_x1_y1,SR_x0_y1,unnamedcast4008USEDMULTIPLEcast,unnamedcast4010USEDMULTIPLEcast,({inp[47:40]}),({inp[39:32]}),({inp[31:24]}),({inp[23:16]}),({inp[15:8]}),({inp[7:0]}),SR_x1_y0,SR_x0_y0};
  // function: process pure=false delay=0
  // function: reset pure=true delay=0
endmodule

module stencilLinebuffer_Auint8_w656_h482_xmin2_ymin2(input CLK, input process_valid, input CE, input [63:0] process_input, output [239:0] process_output, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  wire [191:0] stencilLinebuffer_Auint8_w656_h482_xmin2_ymin2_g_process_output;
  reg process_valid_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay1_validunnamednull0_CECE <= process_valid; end end
  reg process_valid_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay2_validunnamednull0_CECE <= process_valid_delay1_validunnamednull0_CECE; end end
  wire [239:0] stencilLinebuffer_Auint8_w656_h482_xmin2_ymin2_f_process_output;
  assign process_output = stencilLinebuffer_Auint8_w656_h482_xmin2_ymin2_f_process_output;
  // function: process pure=false delay=2
  // function: reset pure=false delay=0
  linebuffer_w656_h482_T8_ymin_2_Auint8 #(.INSTANCE_NAME("stencilLinebuffer_Auint8_w656_h482_xmin2_ymin2_g")) stencilLinebuffer_Auint8_w656_h482_xmin2_ymin2_g(.CLK(CLK), .process_valid(process_valid), .CE(CE), .process_input(process_input), .process_output(stencilLinebuffer_Auint8_w656_h482_xmin2_ymin2_g_process_output), .reset(reset));
  SSR_W3_H3_T8_Auint8 #(.INSTANCE_NAME("stencilLinebuffer_Auint8_w656_h482_xmin2_ymin2_f")) stencilLinebuffer_Auint8_w656_h482_xmin2_ymin2_f(.CLK(CLK), .process_valid(process_valid_delay2_validunnamednull0_CECE), .process_CE(CE), .inp(stencilLinebuffer_Auint8_w656_h482_xmin2_ymin2_g_process_output), .process_output(stencilLinebuffer_Auint8_w656_h482_xmin2_ymin2_f_process_output));
endmodule

module unpackStencil_W3_H3_T8(input CLK, input process_CE, input [239:0] inp, output [575:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [7:0] unnamedcast4522USEDMULTIPLEcast = ({inp[15:8]});
  wire [7:0] unnamedcast4524USEDMULTIPLEcast = ({inp[23:16]});
  wire [7:0] unnamedcast4528USEDMULTIPLEcast = ({inp[95:88]});
  wire [7:0] unnamedcast4530USEDMULTIPLEcast = ({inp[103:96]});
  wire [7:0] unnamedcast4534USEDMULTIPLEcast = ({inp[175:168]});
  wire [7:0] unnamedcast4536USEDMULTIPLEcast = ({inp[183:176]});
  wire [7:0] unnamedcast4542USEDMULTIPLEcast = ({inp[31:24]});
  wire [7:0] unnamedcast4548USEDMULTIPLEcast = ({inp[111:104]});
  wire [7:0] unnamedcast4554USEDMULTIPLEcast = ({inp[191:184]});
  wire [7:0] unnamedcast4560USEDMULTIPLEcast = ({inp[39:32]});
  wire [7:0] unnamedcast4566USEDMULTIPLEcast = ({inp[119:112]});
  wire [7:0] unnamedcast4572USEDMULTIPLEcast = ({inp[199:192]});
  wire [7:0] unnamedcast4578USEDMULTIPLEcast = ({inp[47:40]});
  wire [7:0] unnamedcast4584USEDMULTIPLEcast = ({inp[127:120]});
  wire [7:0] unnamedcast4590USEDMULTIPLEcast = ({inp[207:200]});
  wire [7:0] unnamedcast4596USEDMULTIPLEcast = ({inp[55:48]});
  wire [7:0] unnamedcast4602USEDMULTIPLEcast = ({inp[135:128]});
  wire [7:0] unnamedcast4608USEDMULTIPLEcast = ({inp[215:208]});
  wire [7:0] unnamedcast4614USEDMULTIPLEcast = ({inp[63:56]});
  wire [7:0] unnamedcast4620USEDMULTIPLEcast = ({inp[143:136]});
  wire [7:0] unnamedcast4626USEDMULTIPLEcast = ({inp[223:216]});
  wire [7:0] unnamedcast4632USEDMULTIPLEcast = ({inp[71:64]});
  wire [7:0] unnamedcast4638USEDMULTIPLEcast = ({inp[151:144]});
  wire [7:0] unnamedcast4644USEDMULTIPLEcast = ({inp[231:224]});
  assign process_output = {{({inp[239:232]}),unnamedcast4644USEDMULTIPLEcast,unnamedcast4626USEDMULTIPLEcast,({inp[159:152]}),unnamedcast4638USEDMULTIPLEcast,unnamedcast4620USEDMULTIPLEcast,({inp[79:72]}),unnamedcast4632USEDMULTIPLEcast,unnamedcast4614USEDMULTIPLEcast},{unnamedcast4644USEDMULTIPLEcast,unnamedcast4626USEDMULTIPLEcast,unnamedcast4608USEDMULTIPLEcast,unnamedcast4638USEDMULTIPLEcast,unnamedcast4620USEDMULTIPLEcast,unnamedcast4602USEDMULTIPLEcast,unnamedcast4632USEDMULTIPLEcast,unnamedcast4614USEDMULTIPLEcast,unnamedcast4596USEDMULTIPLEcast},{unnamedcast4626USEDMULTIPLEcast,unnamedcast4608USEDMULTIPLEcast,unnamedcast4590USEDMULTIPLEcast,unnamedcast4620USEDMULTIPLEcast,unnamedcast4602USEDMULTIPLEcast,unnamedcast4584USEDMULTIPLEcast,unnamedcast4614USEDMULTIPLEcast,unnamedcast4596USEDMULTIPLEcast,unnamedcast4578USEDMULTIPLEcast},{unnamedcast4608USEDMULTIPLEcast,unnamedcast4590USEDMULTIPLEcast,unnamedcast4572USEDMULTIPLEcast,unnamedcast4602USEDMULTIPLEcast,unnamedcast4584USEDMULTIPLEcast,unnamedcast4566USEDMULTIPLEcast,unnamedcast4596USEDMULTIPLEcast,unnamedcast4578USEDMULTIPLEcast,unnamedcast4560USEDMULTIPLEcast},{unnamedcast4590USEDMULTIPLEcast,unnamedcast4572USEDMULTIPLEcast,unnamedcast4554USEDMULTIPLEcast,unnamedcast4584USEDMULTIPLEcast,unnamedcast4566USEDMULTIPLEcast,unnamedcast4548USEDMULTIPLEcast,unnamedcast4578USEDMULTIPLEcast,unnamedcast4560USEDMULTIPLEcast,unnamedcast4542USEDMULTIPLEcast},{unnamedcast4572USEDMULTIPLEcast,unnamedcast4554USEDMULTIPLEcast,unnamedcast4536USEDMULTIPLEcast,unnamedcast4566USEDMULTIPLEcast,unnamedcast4548USEDMULTIPLEcast,unnamedcast4530USEDMULTIPLEcast,unnamedcast4560USEDMULTIPLEcast,unnamedcast4542USEDMULTIPLEcast,unnamedcast4524USEDMULTIPLEcast},{unnamedcast4554USEDMULTIPLEcast,unnamedcast4536USEDMULTIPLEcast,unnamedcast4534USEDMULTIPLEcast,unnamedcast4548USEDMULTIPLEcast,unnamedcast4530USEDMULTIPLEcast,unnamedcast4528USEDMULTIPLEcast,unnamedcast4542USEDMULTIPLEcast,unnamedcast4524USEDMULTIPLEcast,unnamedcast4522USEDMULTIPLEcast},{unnamedcast4536USEDMULTIPLEcast,unnamedcast4534USEDMULTIPLEcast,({inp[167:160]}),unnamedcast4530USEDMULTIPLEcast,unnamedcast4528USEDMULTIPLEcast,({inp[87:80]}),unnamedcast4524USEDMULTIPLEcast,unnamedcast4522USEDMULTIPLEcast,({inp[7:0]})}};
  // function: process pure=true delay=0
endmodule

module incif_wrap481_incnil(input CLK, input CE, input [16:0] process_input, output [15:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] unnamedcast3779USEDMULTIPLEcast = (process_input[15:0]);
  assign process_output = (((process_input[16]))?((({(unnamedcast3779USEDMULTIPLEcast==(16'd481))})?((16'd0)):({(unnamedcast3779USEDMULTIPLEcast+(16'd1))}))):(unnamedcast3779USEDMULTIPLEcast));
  // function: process pure=true delay=0
endmodule

module RegBy_incif_wrap481_incnil_CEtrue_init0(input CLK, input set_valid, input CE, input [15:0] set_inp, input setby_valid, input setby_inp, output [15:0] SETBY_OUTPUT, output [15:0] GET_OUTPUT);
parameter INSTANCE_NAME="INST";
  reg [15:0] R = 16'd0;
  wire [15:0] regby_inner_process_output;
  always @(posedge CLK) begin if(set_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(setby_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,set_valid})+({4'b0,setby_valid})) > 5'd1) begin $display("error, function 'set' on instance 'R' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [16:0] unnamedcallArbitrate3830USEDMULTIPLEcallArbitrate = {(set_valid||setby_valid),((set_valid)?(set_inp):(regby_inner_process_output))};
    always @ (posedge CLK) begin if ((unnamedcallArbitrate3830USEDMULTIPLEcallArbitrate[16]) && CE) begin R <= (unnamedcallArbitrate3830USEDMULTIPLEcallArbitrate[15:0]); end end
  assign SETBY_OUTPUT = regby_inner_process_output;
  assign GET_OUTPUT = R;
  // function: set pure=false ONLY WIRE
  // function: setby pure=false ONLY WIRE
  // function: get pure=true ONLY WIRE
  incif_wrap481_incnil #(.INSTANCE_NAME("regby_inner")) regby_inner(.CLK(CLK), .CE(CE), .process_input({setby_inp,R}), .process_output(regby_inner_process_output));
endmodule

module PosSeq_W656_H482_T8(input CLK, input process_valid, input CE, output [255:0] process_output, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  wire [15:0] posX_posSeq_GET_OUTPUT;
  wire [15:0] posY_posSeq_GET_OUTPUT;
  reg [31:0] unnamedtuple3842_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedtuple3842_delay1_validunnamednull0_CECE <= {posY_posSeq_GET_OUTPUT,posX_posSeq_GET_OUTPUT}; end end
  reg [15:0] unnamedbinop3846_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedbinop3846_delay1_validunnamednull0_CECE <= {(posX_posSeq_GET_OUTPUT+(16'd1))}; end end
  reg [15:0] unnamedcall3841_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcall3841_delay1_validunnamednull0_CECE <= posY_posSeq_GET_OUTPUT; end end
  reg [15:0] unnamedbinop3852_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedbinop3852_delay1_validunnamednull0_CECE <= {(posX_posSeq_GET_OUTPUT+(16'd2))}; end end
  reg [15:0] unnamedbinop3858_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedbinop3858_delay1_validunnamednull0_CECE <= {(posX_posSeq_GET_OUTPUT+(16'd3))}; end end
  reg [15:0] unnamedbinop3864_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedbinop3864_delay1_validunnamednull0_CECE <= {(posX_posSeq_GET_OUTPUT+(16'd4))}; end end
  reg [15:0] unnamedbinop3870_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedbinop3870_delay1_validunnamednull0_CECE <= {(posX_posSeq_GET_OUTPUT+(16'd5))}; end end
  reg [15:0] unnamedbinop3876_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedbinop3876_delay1_validunnamednull0_CECE <= {(posX_posSeq_GET_OUTPUT+(16'd6))}; end end
  reg [15:0] unnamedbinop3882_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedbinop3882_delay1_validunnamednull0_CECE <= {(posX_posSeq_GET_OUTPUT+(16'd7))}; end end
  wire [15:0] posX_posSeq_SETBY_OUTPUT;
  wire [15:0] posY_posSeq_SETBY_OUTPUT;
  assign process_output = {{unnamedcall3841_delay1_validunnamednull0_CECE,unnamedbinop3882_delay1_validunnamednull0_CECE},{unnamedcall3841_delay1_validunnamednull0_CECE,unnamedbinop3876_delay1_validunnamednull0_CECE},{unnamedcall3841_delay1_validunnamednull0_CECE,unnamedbinop3870_delay1_validunnamednull0_CECE},{unnamedcall3841_delay1_validunnamednull0_CECE,unnamedbinop3864_delay1_validunnamednull0_CECE},{unnamedcall3841_delay1_validunnamednull0_CECE,unnamedbinop3858_delay1_validunnamednull0_CECE},{unnamedcall3841_delay1_validunnamednull0_CECE,unnamedbinop3852_delay1_validunnamednull0_CECE},{unnamedcall3841_delay1_validunnamednull0_CECE,unnamedbinop3846_delay1_validunnamednull0_CECE},unnamedtuple3842_delay1_validunnamednull0_CECE};
  // function: process pure=false delay=1
  // function: reset pure=false delay=0
  RegBy_incif_wrap648_inc8_CEtrue_init0 #(.INSTANCE_NAME("posX_posSeq")) posX_posSeq(.CLK(CLK), .set_valid(reset), .CE(CE), .set_inp((16'd0)), .setby_valid(process_valid), .setby_inp((1'd1)), .SETBY_OUTPUT(posX_posSeq_SETBY_OUTPUT), .GET_OUTPUT(posX_posSeq_GET_OUTPUT));
  RegBy_incif_wrap481_incnil_CEtrue_init0 #(.INSTANCE_NAME("posY_posSeq")) posY_posSeq(.CLK(CLK), .set_valid(reset), .CE(CE), .set_inp((16'd0)), .setby_valid(process_valid), .setby_inp({(posX_posSeq_GET_OUTPUT==(16'd648))}), .SETBY_OUTPUT(posY_posSeq_SETBY_OUTPUT), .GET_OUTPUT(posY_posSeq_GET_OUTPUT));
endmodule

module packTupleArrays_table__0x42bdcbb0(input CLK, input process_CE, input [831:0] process_input, output [831:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [255:0] unnamedcast3523USEDMULTIPLEcast = (process_input[255:0]);
  wire [575:0] unnamedcast3527USEDMULTIPLEcast = (process_input[831:256]);
  assign process_output = {{({unnamedcast3527USEDMULTIPLEcast[575:504]}),({unnamedcast3523USEDMULTIPLEcast[255:224]})},{({unnamedcast3527USEDMULTIPLEcast[503:432]}),({unnamedcast3523USEDMULTIPLEcast[223:192]})},{({unnamedcast3527USEDMULTIPLEcast[431:360]}),({unnamedcast3523USEDMULTIPLEcast[191:160]})},{({unnamedcast3527USEDMULTIPLEcast[359:288]}),({unnamedcast3523USEDMULTIPLEcast[159:128]})},{({unnamedcast3527USEDMULTIPLEcast[287:216]}),({unnamedcast3523USEDMULTIPLEcast[127:96]})},{({unnamedcast3527USEDMULTIPLEcast[215:144]}),({unnamedcast3523USEDMULTIPLEcast[95:64]})},{({unnamedcast3527USEDMULTIPLEcast[143:72]}),({unnamedcast3523USEDMULTIPLEcast[63:32]})},{({unnamedcast3527USEDMULTIPLEcast[71:0]}),({unnamedcast3523USEDMULTIPLEcast[31:0]})}};
  // function: process pure=true delay=0
endmodule

module index___uint16_uint16__uint8_3_3___1(input CLK, input process_CE, input [103:0] inp, output [71:0] process_output);
parameter INSTANCE_NAME="INST";
  assign process_output = (inp[103:32]);
  // function: process pure=true delay=0
endmodule

module index___uint16_uint16__uint8_3_3___0(input CLK, input process_CE, input [103:0] inp, output [31:0] process_output);
parameter INSTANCE_NAME="INST";
  assign process_output = (inp[31:0]);
  // function: process pure=true delay=0
endmodule

module kern1(input CLK, input process_CE, input [31:0] ksi, output [71:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] unnamedcast2182USEDMULTIPLEcast = (16'd1);
  reg [15:0] unnamedbinop2183_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2183_delay1_validunnamednull0_CEprocess_CE <= {((ksi[15:0])+unnamedcast2182USEDMULTIPLEcast)}; end end
  reg [15:0] unnamedcast2182_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2182_delay1_validunnamednull0_CEprocess_CE <= unnamedcast2182USEDMULTIPLEcast; end end
  reg [15:0] unnamedbinop2186_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2186_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2183_delay1_validunnamednull0_CEprocess_CE&unnamedcast2182_delay1_validunnamednull0_CEprocess_CE)}; end end
  reg [15:0] unnamedbinop2186_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2186_delay2_validunnamednull0_CEprocess_CE <= unnamedbinop2186_delay1_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedbinop2192_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2192_delay1_validunnamednull0_CEprocess_CE <= {((ksi[31:16])+unnamedcast2182USEDMULTIPLEcast)}; end end
  reg [15:0] unnamedbinop2195_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2195_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2192_delay1_validunnamednull0_CEprocess_CE&unnamedcast2182_delay1_validunnamednull0_CEprocess_CE)}; end end
  reg [15:0] unnamedcast2197_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2197_delay1_validunnamednull0_CEprocess_CE <= (16'd2); end end
  reg [15:0] unnamedcast2197_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2197_delay2_validunnamednull0_CEprocess_CE <= unnamedcast2197_delay1_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedbinop2198_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2198_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2195_delay1_validunnamednull0_CEprocess_CE*unnamedcast2197_delay2_validunnamednull0_CEprocess_CE)}; end end
  reg [15:0] unnamedbinop2199_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2199_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2186_delay2_validunnamednull0_CEprocess_CE+unnamedbinop2198_delay1_validunnamednull0_CEprocess_CE)}; end end
  reg [15:0] unnamedcast2205_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2205_delay1_validunnamednull0_CEprocess_CE <= (16'd0); end end
  reg [15:0] unnamedcast2205_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2205_delay2_validunnamednull0_CEprocess_CE <= unnamedcast2205_delay1_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedcast2205_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2205_delay3_validunnamednull0_CEprocess_CE <= unnamedcast2205_delay2_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedcast2205_delay4_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2205_delay4_validunnamednull0_CEprocess_CE <= unnamedcast2205_delay3_validunnamednull0_CEprocess_CE; end end
  reg unnamedbinop2206_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2206_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2199_delay1_validunnamednull0_CEprocess_CE==unnamedcast2205_delay4_validunnamednull0_CEprocess_CE)}; end end
  wire [72:0] unnamedtuple2207USEDMULTIPLEtuple = {unnamedbinop2206_delay1_validunnamednull0_CEprocess_CE,({8'd0, 8'd0, 8'd0, 8'd2, 8'd0, 8'd2, 8'd0, 8'd0, 8'd0})};
  reg [15:0] unnamedcast2182_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2182_delay2_validunnamednull0_CEprocess_CE <= unnamedcast2182_delay1_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedcast2182_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2182_delay3_validunnamednull0_CEprocess_CE <= unnamedcast2182_delay2_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedcast2182_delay4_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2182_delay4_validunnamednull0_CEprocess_CE <= unnamedcast2182_delay3_validunnamednull0_CEprocess_CE; end end
  reg unnamedbinop2210_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2210_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2199_delay1_validunnamednull0_CEprocess_CE==unnamedcast2182_delay4_validunnamednull0_CEprocess_CE)}; end end
  reg [72:0] unnamedselect2222_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedselect2222_delay1_validunnamednull0_CEprocess_CE <= (((unnamedtuple2207USEDMULTIPLEtuple[72]))?(unnamedtuple2207USEDMULTIPLEtuple):({unnamedbinop2210_delay1_validunnamednull0_CEprocess_CE,({8'd0, 8'd0, 8'd0, 8'd0, 8'd4, 8'd0, 8'd0, 8'd0, 8'd0})})); end end
  reg [15:0] unnamedcast2197_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2197_delay3_validunnamednull0_CEprocess_CE <= unnamedcast2197_delay2_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedcast2197_delay4_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2197_delay4_validunnamednull0_CEprocess_CE <= unnamedcast2197_delay3_validunnamednull0_CEprocess_CE; end end
  reg unnamedbinop2214_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2214_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2199_delay1_validunnamednull0_CEprocess_CE==unnamedcast2197_delay4_validunnamednull0_CEprocess_CE)}; end end
  wire [72:0] unnamedtuple2215USEDMULTIPLEtuple = {unnamedbinop2214_delay1_validunnamednull0_CEprocess_CE,({8'd1, 8'd0, 8'd1, 8'd0, 8'd0, 8'd0, 8'd1, 8'd0, 8'd1})};
  reg [15:0] unnamedcast2217_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2217_delay1_validunnamednull0_CEprocess_CE <= (16'd3); end end
  reg [15:0] unnamedcast2217_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2217_delay2_validunnamednull0_CEprocess_CE <= unnamedcast2217_delay1_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedcast2217_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2217_delay3_validunnamednull0_CEprocess_CE <= unnamedcast2217_delay2_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedcast2217_delay4_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2217_delay4_validunnamednull0_CEprocess_CE <= unnamedcast2217_delay3_validunnamednull0_CEprocess_CE; end end
  reg unnamedbinop2218_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2218_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2199_delay1_validunnamednull0_CEprocess_CE==unnamedcast2217_delay4_validunnamednull0_CEprocess_CE)}; end end
  reg [72:0] unnamedselect2225_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedselect2225_delay1_validunnamednull0_CEprocess_CE <= (((unnamedtuple2215USEDMULTIPLEtuple[72]))?(unnamedtuple2215USEDMULTIPLEtuple):({unnamedbinop2218_delay1_validunnamednull0_CEprocess_CE,({8'd0, 8'd2, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd2, 8'd0})})); end end
  reg [72:0] unnamedselect2228_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedselect2228_delay1_validunnamednull0_CEprocess_CE <= (((unnamedselect2222_delay1_validunnamednull0_CEprocess_CE[72]))?(unnamedselect2222_delay1_validunnamednull0_CEprocess_CE):(unnamedselect2225_delay1_validunnamednull0_CEprocess_CE)); end end
  assign process_output = (unnamedselect2228_delay1_validunnamednull0_CEprocess_CE[71:0]);
  // function: process pure=true delay=7
endmodule

module packTupleArrays_table__0x410fe0f0(input CLK, input process_CE, input [143:0] process_input, output [143:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [71:0] unnamedcast2325USEDMULTIPLEcast = (process_input[71:0]);
  wire [71:0] unnamedcast2329USEDMULTIPLEcast = (process_input[143:72]);
  assign process_output = {{({unnamedcast2329USEDMULTIPLEcast[71:64]}),({unnamedcast2325USEDMULTIPLEcast[71:64]})},{({unnamedcast2329USEDMULTIPLEcast[63:56]}),({unnamedcast2325USEDMULTIPLEcast[63:56]})},{({unnamedcast2329USEDMULTIPLEcast[55:48]}),({unnamedcast2325USEDMULTIPLEcast[55:48]})},{({unnamedcast2329USEDMULTIPLEcast[47:40]}),({unnamedcast2325USEDMULTIPLEcast[47:40]})},{({unnamedcast2329USEDMULTIPLEcast[39:32]}),({unnamedcast2325USEDMULTIPLEcast[39:32]})},{({unnamedcast2329USEDMULTIPLEcast[31:24]}),({unnamedcast2325USEDMULTIPLEcast[31:24]})},{({unnamedcast2329USEDMULTIPLEcast[23:16]}),({unnamedcast2325USEDMULTIPLEcast[23:16]})},{({unnamedcast2329USEDMULTIPLEcast[15:8]}),({unnamedcast2325USEDMULTIPLEcast[15:8]})},{({unnamedcast2329USEDMULTIPLEcast[7:0]}),({unnamedcast2325USEDMULTIPLEcast[7:0]})}};
  // function: process pure=true delay=0
endmodule

module partial_mult(input CLK, input process_CE, input [15:0] inp, output [15:0] process_output);
parameter INSTANCE_NAME="INST";
  reg [15:0] unnamedbinop2413_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2413_delay1_validunnamednull0_CEprocess_CE <= {({8'b0,(inp[7:0])}*{8'b0,(inp[15:8])})}; end end
  assign process_output = unnamedbinop2413_delay1_validunnamednull0_CEprocess_CE;
  // function: process pure=true delay=1
endmodule

module map_partial_mult_W3_H3(input CLK, input process_CE, input [143:0] process_input, output [143:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] inner0_0_process_output;
  wire [15:0] inner1_0_process_output;
  wire [15:0] inner2_0_process_output;
  wire [15:0] inner0_1_process_output;
  wire [15:0] inner1_1_process_output;
  wire [15:0] inner2_1_process_output;
  wire [15:0] inner0_2_process_output;
  wire [15:0] inner1_2_process_output;
  wire [15:0] inner2_2_process_output;
  assign process_output = {inner2_2_process_output,inner1_2_process_output,inner0_2_process_output,inner2_1_process_output,inner1_1_process_output,inner0_1_process_output,inner2_0_process_output,inner1_0_process_output,inner0_0_process_output};
  // function: process pure=true delay=1
  partial_mult #(.INSTANCE_NAME("inner0_0")) inner0_0(.CLK(CLK), .process_CE(process_CE), .inp(({process_input[15:0]})), .process_output(inner0_0_process_output));
  partial_mult #(.INSTANCE_NAME("inner1_0")) inner1_0(.CLK(CLK), .process_CE(process_CE), .inp(({process_input[31:16]})), .process_output(inner1_0_process_output));
  partial_mult #(.INSTANCE_NAME("inner2_0")) inner2_0(.CLK(CLK), .process_CE(process_CE), .inp(({process_input[47:32]})), .process_output(inner2_0_process_output));
  partial_mult #(.INSTANCE_NAME("inner0_1")) inner0_1(.CLK(CLK), .process_CE(process_CE), .inp(({process_input[63:48]})), .process_output(inner0_1_process_output));
  partial_mult #(.INSTANCE_NAME("inner1_1")) inner1_1(.CLK(CLK), .process_CE(process_CE), .inp(({process_input[79:64]})), .process_output(inner1_1_process_output));
  partial_mult #(.INSTANCE_NAME("inner2_1")) inner2_1(.CLK(CLK), .process_CE(process_CE), .inp(({process_input[95:80]})), .process_output(inner2_1_process_output));
  partial_mult #(.INSTANCE_NAME("inner0_2")) inner0_2(.CLK(CLK), .process_CE(process_CE), .inp(({process_input[111:96]})), .process_output(inner0_2_process_output));
  partial_mult #(.INSTANCE_NAME("inner1_2")) inner1_2(.CLK(CLK), .process_CE(process_CE), .inp(({process_input[127:112]})), .process_output(inner1_2_process_output));
  partial_mult #(.INSTANCE_NAME("inner2_2")) inner2_2(.CLK(CLK), .process_CE(process_CE), .inp(({process_input[143:128]})), .process_output(inner2_2_process_output));
endmodule

module sum(input CLK, input process_CE, input [31:0] inp, output [15:0] process_output);
parameter INSTANCE_NAME="INST";
  reg [15:0] unnamedbinop2461_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2461_delay1_validunnamednull0_CEprocess_CE <= {((inp[15:0])+(inp[31:16]))}; end end
  assign process_output = unnamedbinop2461_delay1_validunnamednull0_CEprocess_CE;
  // function: process pure=true delay=1
endmodule

module reduce_sum_W3_H3(input CLK, input process_CE, input [143:0] process_input, output [15:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] inner0_process_output;
  wire [15:0] inner1_process_output;
  wire [15:0] inner4_process_output;
  wire [15:0] inner2_process_output;
  wire [15:0] inner3_process_output;
  wire [15:0] inner5_process_output;
  wire [15:0] inner6_process_output;
  reg [15:0] unnamedcast2491_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2491_delay1_validunnamednull0_CEprocess_CE <= ({process_input[143:128]}); end end
  reg [15:0] unnamedcast2491_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2491_delay2_validunnamednull0_CEprocess_CE <= unnamedcast2491_delay1_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedcast2491_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2491_delay3_validunnamednull0_CEprocess_CE <= unnamedcast2491_delay2_validunnamednull0_CEprocess_CE; end end
  wire [15:0] inner7_process_output;
  assign process_output = inner7_process_output;
  // function: process pure=true delay=4
  sum #(.INSTANCE_NAME("inner0")) inner0(.CLK(CLK), .process_CE(process_CE), .inp({({process_input[31:16]}),({process_input[15:0]})}), .process_output(inner0_process_output));
  sum #(.INSTANCE_NAME("inner1")) inner1(.CLK(CLK), .process_CE(process_CE), .inp({({process_input[63:48]}),({process_input[47:32]})}), .process_output(inner1_process_output));
  sum #(.INSTANCE_NAME("inner2")) inner2(.CLK(CLK), .process_CE(process_CE), .inp({({process_input[95:80]}),({process_input[79:64]})}), .process_output(inner2_process_output));
  sum #(.INSTANCE_NAME("inner3")) inner3(.CLK(CLK), .process_CE(process_CE), .inp({({process_input[127:112]}),({process_input[111:96]})}), .process_output(inner3_process_output));
  sum #(.INSTANCE_NAME("inner4")) inner4(.CLK(CLK), .process_CE(process_CE), .inp({inner1_process_output,inner0_process_output}), .process_output(inner4_process_output));
  sum #(.INSTANCE_NAME("inner5")) inner5(.CLK(CLK), .process_CE(process_CE), .inp({inner3_process_output,inner2_process_output}), .process_output(inner5_process_output));
  sum #(.INSTANCE_NAME("inner6")) inner6(.CLK(CLK), .process_CE(process_CE), .inp({inner5_process_output,inner4_process_output}), .process_output(inner6_process_output));
  sum #(.INSTANCE_NAME("inner7")) inner7(.CLK(CLK), .process_CE(process_CE), .inp({unnamedcast2491_delay3_validunnamednull0_CEprocess_CE,inner6_process_output}), .process_output(inner7_process_output));
endmodule

module touint8(input CLK, input process_CE, input [15:0] inp, output [7:0] process_output);
parameter INSTANCE_NAME="INST";
  reg [15:0] unnamedbinop2510_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2510_delay1_validunnamednull0_CEprocess_CE <= {(inp>>>(16'd2))}; end end
  reg [15:0] unnamedcast2512_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2512_delay1_validunnamednull0_CEprocess_CE <= (16'd255); end end
  reg unnamedbinop2513_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2513_delay1_validunnamednull0_CEprocess_CE <= {((unnamedbinop2510_delay1_validunnamednull0_CEprocess_CE)>(unnamedcast2512_delay1_validunnamednull0_CEprocess_CE))}; end end
  reg [7:0] unnamedcast2516_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2516_delay1_validunnamednull0_CEprocess_CE <= (8'd255); end end
  reg [7:0] unnamedcast2516_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2516_delay2_validunnamednull0_CEprocess_CE <= unnamedcast2516_delay1_validunnamednull0_CEprocess_CE; end end
  reg [7:0] unnamedcast2515_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2515_delay1_validunnamednull0_CEprocess_CE <= unnamedbinop2510_delay1_validunnamednull0_CEprocess_CE[7:0]; end end
  reg [7:0] unnamedselect2517_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedselect2517_delay1_validunnamednull0_CEprocess_CE <= ((unnamedbinop2513_delay1_validunnamednull0_CEprocess_CE)?(unnamedcast2516_delay2_validunnamednull0_CEprocess_CE):(unnamedcast2515_delay1_validunnamednull0_CEprocess_CE)); end end
  assign process_output = unnamedselect2517_delay1_validunnamednull0_CEprocess_CE;
  // function: process pure=true delay=3
endmodule

module kern2(input CLK, input process_CE, input [31:0] ksi, output [71:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] unnamedcast2543USEDMULTIPLEcast = (16'd1);
  reg [15:0] unnamedbinop2544_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2544_delay1_validunnamednull0_CEprocess_CE <= {((ksi[15:0])+unnamedcast2543USEDMULTIPLEcast)}; end end
  reg [15:0] unnamedcast2543_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2543_delay1_validunnamednull0_CEprocess_CE <= unnamedcast2543USEDMULTIPLEcast; end end
  reg [15:0] unnamedbinop2547_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2547_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2544_delay1_validunnamednull0_CEprocess_CE&unnamedcast2543_delay1_validunnamednull0_CEprocess_CE)}; end end
  reg [15:0] unnamedbinop2547_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2547_delay2_validunnamednull0_CEprocess_CE <= unnamedbinop2547_delay1_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedbinop2553_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2553_delay1_validunnamednull0_CEprocess_CE <= {((ksi[31:16])+unnamedcast2543USEDMULTIPLEcast)}; end end
  reg [15:0] unnamedbinop2556_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2556_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2553_delay1_validunnamednull0_CEprocess_CE&unnamedcast2543_delay1_validunnamednull0_CEprocess_CE)}; end end
  reg [15:0] unnamedcast2558_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2558_delay1_validunnamednull0_CEprocess_CE <= (16'd2); end end
  reg [15:0] unnamedcast2558_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2558_delay2_validunnamednull0_CEprocess_CE <= unnamedcast2558_delay1_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedbinop2559_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2559_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2556_delay1_validunnamednull0_CEprocess_CE*unnamedcast2558_delay2_validunnamednull0_CEprocess_CE)}; end end
  reg [15:0] unnamedbinop2560_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2560_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2547_delay2_validunnamednull0_CEprocess_CE+unnamedbinop2559_delay1_validunnamednull0_CEprocess_CE)}; end end
  reg [15:0] unnamedcast2566_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2566_delay1_validunnamednull0_CEprocess_CE <= (16'd0); end end
  reg [15:0] unnamedcast2566_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2566_delay2_validunnamednull0_CEprocess_CE <= unnamedcast2566_delay1_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedcast2566_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2566_delay3_validunnamednull0_CEprocess_CE <= unnamedcast2566_delay2_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedcast2566_delay4_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2566_delay4_validunnamednull0_CEprocess_CE <= unnamedcast2566_delay3_validunnamednull0_CEprocess_CE; end end
  reg unnamedbinop2567_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2567_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2560_delay1_validunnamednull0_CEprocess_CE==unnamedcast2566_delay4_validunnamednull0_CEprocess_CE)}; end end
  wire [72:0] unnamedtuple2568USEDMULTIPLEtuple = {unnamedbinop2567_delay1_validunnamednull0_CEprocess_CE,({8'd0, 8'd0, 8'd0, 8'd0, 8'd4, 8'd0, 8'd0, 8'd0, 8'd0})};
  reg [15:0] unnamedcast2543_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2543_delay2_validunnamednull0_CEprocess_CE <= unnamedcast2543_delay1_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedcast2543_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2543_delay3_validunnamednull0_CEprocess_CE <= unnamedcast2543_delay2_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedcast2543_delay4_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2543_delay4_validunnamednull0_CEprocess_CE <= unnamedcast2543_delay3_validunnamednull0_CEprocess_CE; end end
  reg unnamedbinop2571_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2571_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2560_delay1_validunnamednull0_CEprocess_CE==unnamedcast2543_delay4_validunnamednull0_CEprocess_CE)}; end end
  reg [72:0] unnamedselect2583_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedselect2583_delay1_validunnamednull0_CEprocess_CE <= (((unnamedtuple2568USEDMULTIPLEtuple[72]))?(unnamedtuple2568USEDMULTIPLEtuple):({unnamedbinop2571_delay1_validunnamednull0_CEprocess_CE,({8'd0, 8'd1, 8'd0, 8'd1, 8'd0, 8'd1, 8'd0, 8'd1, 8'd0})})); end end
  reg [15:0] unnamedcast2558_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2558_delay3_validunnamednull0_CEprocess_CE <= unnamedcast2558_delay2_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedcast2558_delay4_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2558_delay4_validunnamednull0_CEprocess_CE <= unnamedcast2558_delay3_validunnamednull0_CEprocess_CE; end end
  reg unnamedbinop2575_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2575_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2560_delay1_validunnamednull0_CEprocess_CE==unnamedcast2558_delay4_validunnamednull0_CEprocess_CE)}; end end
  wire [72:0] unnamedtuple2576USEDMULTIPLEtuple = {unnamedbinop2575_delay1_validunnamednull0_CEprocess_CE,({8'd0, 8'd1, 8'd0, 8'd1, 8'd0, 8'd1, 8'd0, 8'd1, 8'd0})};
  reg [15:0] unnamedcast2578_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2578_delay1_validunnamednull0_CEprocess_CE <= (16'd3); end end
  reg [15:0] unnamedcast2578_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2578_delay2_validunnamednull0_CEprocess_CE <= unnamedcast2578_delay1_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedcast2578_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2578_delay3_validunnamednull0_CEprocess_CE <= unnamedcast2578_delay2_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedcast2578_delay4_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2578_delay4_validunnamednull0_CEprocess_CE <= unnamedcast2578_delay3_validunnamednull0_CEprocess_CE; end end
  reg unnamedbinop2579_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2579_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2560_delay1_validunnamednull0_CEprocess_CE==unnamedcast2578_delay4_validunnamednull0_CEprocess_CE)}; end end
  reg [72:0] unnamedselect2586_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedselect2586_delay1_validunnamednull0_CEprocess_CE <= (((unnamedtuple2576USEDMULTIPLEtuple[72]))?(unnamedtuple2576USEDMULTIPLEtuple):({unnamedbinop2579_delay1_validunnamednull0_CEprocess_CE,({8'd0, 8'd0, 8'd0, 8'd0, 8'd4, 8'd0, 8'd0, 8'd0, 8'd0})})); end end
  reg [72:0] unnamedselect2589_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedselect2589_delay1_validunnamednull0_CEprocess_CE <= (((unnamedselect2583_delay1_validunnamednull0_CEprocess_CE[72]))?(unnamedselect2583_delay1_validunnamednull0_CEprocess_CE):(unnamedselect2586_delay1_validunnamednull0_CEprocess_CE)); end end
  assign process_output = (unnamedselect2589_delay1_validunnamednull0_CEprocess_CE[71:0]);
  // function: process pure=true delay=7
endmodule

module packTupleArrays_table__0x423f0260(input CLK, input process_CE, input [143:0] process_input, output [143:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [71:0] unnamedcast2686USEDMULTIPLEcast = (process_input[71:0]);
  wire [71:0] unnamedcast2690USEDMULTIPLEcast = (process_input[143:72]);
  assign process_output = {{({unnamedcast2690USEDMULTIPLEcast[71:64]}),({unnamedcast2686USEDMULTIPLEcast[71:64]})},{({unnamedcast2690USEDMULTIPLEcast[63:56]}),({unnamedcast2686USEDMULTIPLEcast[63:56]})},{({unnamedcast2690USEDMULTIPLEcast[55:48]}),({unnamedcast2686USEDMULTIPLEcast[55:48]})},{({unnamedcast2690USEDMULTIPLEcast[47:40]}),({unnamedcast2686USEDMULTIPLEcast[47:40]})},{({unnamedcast2690USEDMULTIPLEcast[39:32]}),({unnamedcast2686USEDMULTIPLEcast[39:32]})},{({unnamedcast2690USEDMULTIPLEcast[31:24]}),({unnamedcast2686USEDMULTIPLEcast[31:24]})},{({unnamedcast2690USEDMULTIPLEcast[23:16]}),({unnamedcast2686USEDMULTIPLEcast[23:16]})},{({unnamedcast2690USEDMULTIPLEcast[15:8]}),({unnamedcast2686USEDMULTIPLEcast[15:8]})},{({unnamedcast2690USEDMULTIPLEcast[7:0]}),({unnamedcast2686USEDMULTIPLEcast[7:0]})}};
  // function: process pure=true delay=0
endmodule

module kern3(input CLK, input process_CE, input [31:0] ksi, output [71:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] unnamedcast2772USEDMULTIPLEcast = (16'd1);
  reg [15:0] unnamedbinop2773_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2773_delay1_validunnamednull0_CEprocess_CE <= {((ksi[15:0])+unnamedcast2772USEDMULTIPLEcast)}; end end
  reg [15:0] unnamedcast2772_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2772_delay1_validunnamednull0_CEprocess_CE <= unnamedcast2772USEDMULTIPLEcast; end end
  reg [15:0] unnamedbinop2776_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2776_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2773_delay1_validunnamednull0_CEprocess_CE&unnamedcast2772_delay1_validunnamednull0_CEprocess_CE)}; end end
  reg [15:0] unnamedbinop2776_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2776_delay2_validunnamednull0_CEprocess_CE <= unnamedbinop2776_delay1_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedbinop2782_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2782_delay1_validunnamednull0_CEprocess_CE <= {((ksi[31:16])+unnamedcast2772USEDMULTIPLEcast)}; end end
  reg [15:0] unnamedbinop2785_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2785_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2782_delay1_validunnamednull0_CEprocess_CE&unnamedcast2772_delay1_validunnamednull0_CEprocess_CE)}; end end
  reg [15:0] unnamedcast2787_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2787_delay1_validunnamednull0_CEprocess_CE <= (16'd2); end end
  reg [15:0] unnamedcast2787_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2787_delay2_validunnamednull0_CEprocess_CE <= unnamedcast2787_delay1_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedbinop2788_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2788_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2785_delay1_validunnamednull0_CEprocess_CE*unnamedcast2787_delay2_validunnamednull0_CEprocess_CE)}; end end
  reg [15:0] unnamedbinop2789_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2789_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2776_delay2_validunnamednull0_CEprocess_CE+unnamedbinop2788_delay1_validunnamednull0_CEprocess_CE)}; end end
  reg [15:0] unnamedcast2795_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2795_delay1_validunnamednull0_CEprocess_CE <= (16'd0); end end
  reg [15:0] unnamedcast2795_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2795_delay2_validunnamednull0_CEprocess_CE <= unnamedcast2795_delay1_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedcast2795_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2795_delay3_validunnamednull0_CEprocess_CE <= unnamedcast2795_delay2_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedcast2795_delay4_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2795_delay4_validunnamednull0_CEprocess_CE <= unnamedcast2795_delay3_validunnamednull0_CEprocess_CE; end end
  reg unnamedbinop2796_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2796_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2789_delay1_validunnamednull0_CEprocess_CE==unnamedcast2795_delay4_validunnamednull0_CEprocess_CE)}; end end
  wire [72:0] unnamedtuple2797USEDMULTIPLEtuple = {unnamedbinop2796_delay1_validunnamednull0_CEprocess_CE,({8'd0, 8'd2, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd2, 8'd0})};
  reg [15:0] unnamedcast2772_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2772_delay2_validunnamednull0_CEprocess_CE <= unnamedcast2772_delay1_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedcast2772_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2772_delay3_validunnamednull0_CEprocess_CE <= unnamedcast2772_delay2_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedcast2772_delay4_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2772_delay4_validunnamednull0_CEprocess_CE <= unnamedcast2772_delay3_validunnamednull0_CEprocess_CE; end end
  reg unnamedbinop2800_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2800_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2789_delay1_validunnamednull0_CEprocess_CE==unnamedcast2772_delay4_validunnamednull0_CEprocess_CE)}; end end
  reg [72:0] unnamedselect2812_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedselect2812_delay1_validunnamednull0_CEprocess_CE <= (((unnamedtuple2797USEDMULTIPLEtuple[72]))?(unnamedtuple2797USEDMULTIPLEtuple):({unnamedbinop2800_delay1_validunnamednull0_CEprocess_CE,({8'd1, 8'd0, 8'd1, 8'd0, 8'd0, 8'd0, 8'd1, 8'd0, 8'd1})})); end end
  reg [15:0] unnamedcast2787_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2787_delay3_validunnamednull0_CEprocess_CE <= unnamedcast2787_delay2_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedcast2787_delay4_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2787_delay4_validunnamednull0_CEprocess_CE <= unnamedcast2787_delay3_validunnamednull0_CEprocess_CE; end end
  reg unnamedbinop2804_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2804_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2789_delay1_validunnamednull0_CEprocess_CE==unnamedcast2787_delay4_validunnamednull0_CEprocess_CE)}; end end
  wire [72:0] unnamedtuple2805USEDMULTIPLEtuple = {unnamedbinop2804_delay1_validunnamednull0_CEprocess_CE,({8'd0, 8'd0, 8'd0, 8'd0, 8'd4, 8'd0, 8'd0, 8'd0, 8'd0})};
  reg [15:0] unnamedcast2807_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2807_delay1_validunnamednull0_CEprocess_CE <= (16'd3); end end
  reg [15:0] unnamedcast2807_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2807_delay2_validunnamednull0_CEprocess_CE <= unnamedcast2807_delay1_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedcast2807_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2807_delay3_validunnamednull0_CEprocess_CE <= unnamedcast2807_delay2_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedcast2807_delay4_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast2807_delay4_validunnamednull0_CEprocess_CE <= unnamedcast2807_delay3_validunnamednull0_CEprocess_CE; end end
  reg unnamedbinop2808_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop2808_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop2789_delay1_validunnamednull0_CEprocess_CE==unnamedcast2807_delay4_validunnamednull0_CEprocess_CE)}; end end
  reg [72:0] unnamedselect2815_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedselect2815_delay1_validunnamednull0_CEprocess_CE <= (((unnamedtuple2805USEDMULTIPLEtuple[72]))?(unnamedtuple2805USEDMULTIPLEtuple):({unnamedbinop2808_delay1_validunnamednull0_CEprocess_CE,({8'd0, 8'd0, 8'd0, 8'd2, 8'd0, 8'd2, 8'd0, 8'd0, 8'd0})})); end end
  reg [72:0] unnamedselect2818_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedselect2818_delay1_validunnamednull0_CEprocess_CE <= (((unnamedselect2812_delay1_validunnamednull0_CEprocess_CE[72]))?(unnamedselect2812_delay1_validunnamednull0_CEprocess_CE):(unnamedselect2815_delay1_validunnamednull0_CEprocess_CE)); end end
  assign process_output = (unnamedselect2818_delay1_validunnamednull0_CEprocess_CE[71:0]);
  // function: process pure=true delay=7
endmodule

module packTupleArrays_table__0x42d99dd8(input CLK, input process_CE, input [143:0] process_input, output [143:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [71:0] unnamedcast2915USEDMULTIPLEcast = (process_input[71:0]);
  wire [71:0] unnamedcast2919USEDMULTIPLEcast = (process_input[143:72]);
  assign process_output = {{({unnamedcast2919USEDMULTIPLEcast[71:64]}),({unnamedcast2915USEDMULTIPLEcast[71:64]})},{({unnamedcast2919USEDMULTIPLEcast[63:56]}),({unnamedcast2915USEDMULTIPLEcast[63:56]})},{({unnamedcast2919USEDMULTIPLEcast[55:48]}),({unnamedcast2915USEDMULTIPLEcast[55:48]})},{({unnamedcast2919USEDMULTIPLEcast[47:40]}),({unnamedcast2915USEDMULTIPLEcast[47:40]})},{({unnamedcast2919USEDMULTIPLEcast[39:32]}),({unnamedcast2915USEDMULTIPLEcast[39:32]})},{({unnamedcast2919USEDMULTIPLEcast[31:24]}),({unnamedcast2915USEDMULTIPLEcast[31:24]})},{({unnamedcast2919USEDMULTIPLEcast[23:16]}),({unnamedcast2915USEDMULTIPLEcast[23:16]})},{({unnamedcast2919USEDMULTIPLEcast[15:8]}),({unnamedcast2915USEDMULTIPLEcast[15:8]})},{({unnamedcast2919USEDMULTIPLEcast[7:0]}),({unnamedcast2915USEDMULTIPLEcast[7:0]})}};
  // function: process pure=true delay=0
endmodule

module dem(input CLK, input CE, input [103:0] process_input, output [23:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [71:0] dat_process_output;
  reg [71:0] unnamedcall2997_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcall2997_delay1_validunnamednull0_CECE <= dat_process_output; end end
  reg [71:0] unnamedcall2997_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcall2997_delay2_validunnamednull0_CECE <= unnamedcall2997_delay1_validunnamednull0_CECE; end end
  reg [71:0] unnamedcall2997_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcall2997_delay3_validunnamednull0_CECE <= unnamedcall2997_delay2_validunnamednull0_CECE; end end
  reg [71:0] unnamedcall2997_delay4_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcall2997_delay4_validunnamednull0_CECE <= unnamedcall2997_delay3_validunnamednull0_CECE; end end
  reg [71:0] unnamedcall2997_delay5_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcall2997_delay5_validunnamednull0_CECE <= unnamedcall2997_delay4_validunnamednull0_CECE; end end
  reg [71:0] unnamedcall2997_delay6_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcall2997_delay6_validunnamednull0_CECE <= unnamedcall2997_delay5_validunnamednull0_CECE; end end
  reg [71:0] unnamedcall2997_delay7_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcall2997_delay7_validunnamednull0_CECE <= unnamedcall2997_delay6_validunnamednull0_CECE; end end
  wire [31:0] xy_process_output;
  wire [71:0] k1_process_output;
  wire [143:0] packedtup1_process_output;
  wire [143:0] partialll1_process_output;
  wire [15:0] sum1_process_output;
  wire [7:0] touint81_process_output;
  wire [71:0] k2_process_output;
  wire [143:0] packedtup2_process_output;
  wire [143:0] partialll2_process_output;
  wire [15:0] sum2_process_output;
  wire [7:0] touint82_process_output;
  wire [71:0] k3_process_output;
  wire [143:0] packedtup3_process_output;
  wire [143:0] partialll3_process_output;
  wire [15:0] sum3_process_output;
  wire [7:0] touint83_process_output;
  assign process_output = {touint83_process_output,touint82_process_output,touint81_process_output};
  // function: process pure=true delay=15
  // function: reset pure=true delay=0
  index___uint16_uint16__uint8_3_3___1 #(.INSTANCE_NAME("dat")) dat(.CLK(CLK), .process_CE(CE), .inp(process_input), .process_output(dat_process_output));
  index___uint16_uint16__uint8_3_3___0 #(.INSTANCE_NAME("xy")) xy(.CLK(CLK), .process_CE(CE), .inp(process_input), .process_output(xy_process_output));
  kern1 #(.INSTANCE_NAME("k1")) k1(.CLK(CLK), .process_CE(CE), .ksi(xy_process_output), .process_output(k1_process_output));
  packTupleArrays_table__0x410fe0f0 #(.INSTANCE_NAME("packedtup1")) packedtup1(.CLK(CLK), .process_CE(CE), .process_input({k1_process_output,unnamedcall2997_delay7_validunnamednull0_CECE}), .process_output(packedtup1_process_output));
  map_partial_mult_W3_H3 #(.INSTANCE_NAME("partialll1")) partialll1(.CLK(CLK), .process_CE(CE), .process_input(packedtup1_process_output), .process_output(partialll1_process_output));
  reduce_sum_W3_H3 #(.INSTANCE_NAME("sum1")) sum1(.CLK(CLK), .process_CE(CE), .process_input(partialll1_process_output), .process_output(sum1_process_output));
  touint8 #(.INSTANCE_NAME("touint81")) touint81(.CLK(CLK), .process_CE(CE), .inp(sum1_process_output), .process_output(touint81_process_output));
  kern2 #(.INSTANCE_NAME("k2")) k2(.CLK(CLK), .process_CE(CE), .ksi(xy_process_output), .process_output(k2_process_output));
  packTupleArrays_table__0x423f0260 #(.INSTANCE_NAME("packedtup2")) packedtup2(.CLK(CLK), .process_CE(CE), .process_input({k2_process_output,unnamedcall2997_delay7_validunnamednull0_CECE}), .process_output(packedtup2_process_output));
  map_partial_mult_W3_H3 #(.INSTANCE_NAME("partialll2")) partialll2(.CLK(CLK), .process_CE(CE), .process_input(packedtup2_process_output), .process_output(partialll2_process_output));
  reduce_sum_W3_H3 #(.INSTANCE_NAME("sum2")) sum2(.CLK(CLK), .process_CE(CE), .process_input(partialll2_process_output), .process_output(sum2_process_output));
  touint8 #(.INSTANCE_NAME("touint82")) touint82(.CLK(CLK), .process_CE(CE), .inp(sum2_process_output), .process_output(touint82_process_output));
  kern3 #(.INSTANCE_NAME("k3")) k3(.CLK(CLK), .process_CE(CE), .ksi(xy_process_output), .process_output(k3_process_output));
  packTupleArrays_table__0x42d99dd8 #(.INSTANCE_NAME("packedtup3")) packedtup3(.CLK(CLK), .process_CE(CE), .process_input({k3_process_output,unnamedcall2997_delay7_validunnamednull0_CECE}), .process_output(packedtup3_process_output));
  map_partial_mult_W3_H3 #(.INSTANCE_NAME("partialll3")) partialll3(.CLK(CLK), .process_CE(CE), .process_input(packedtup3_process_output), .process_output(partialll3_process_output));
  reduce_sum_W3_H3 #(.INSTANCE_NAME("sum3")) sum3(.CLK(CLK), .process_CE(CE), .process_input(partialll3_process_output), .process_output(sum3_process_output));
  touint8 #(.INSTANCE_NAME("touint83")) touint83(.CLK(CLK), .process_CE(CE), .inp(sum3_process_output), .process_output(touint83_process_output));
endmodule

module map_dem_W8_H1(input CLK, input process_CE, input [831:0] process_input, output [191:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [23:0] inner0_0_process_output;
  wire [23:0] inner1_0_process_output;
  wire [23:0] inner2_0_process_output;
  wire [23:0] inner3_0_process_output;
  wire [23:0] inner4_0_process_output;
  wire [23:0] inner5_0_process_output;
  wire [23:0] inner6_0_process_output;
  wire [23:0] inner7_0_process_output;
  assign process_output = {inner7_0_process_output,inner6_0_process_output,inner5_0_process_output,inner4_0_process_output,inner3_0_process_output,inner2_0_process_output,inner1_0_process_output,inner0_0_process_output};
  // function: process pure=true delay=15
  dem #(.INSTANCE_NAME("inner0_0")) inner0_0(.CLK(CLK), .CE(process_CE), .process_input(({process_input[103:0]})), .process_output(inner0_0_process_output));
  dem #(.INSTANCE_NAME("inner1_0")) inner1_0(.CLK(CLK), .CE(process_CE), .process_input(({process_input[207:104]})), .process_output(inner1_0_process_output));
  dem #(.INSTANCE_NAME("inner2_0")) inner2_0(.CLK(CLK), .CE(process_CE), .process_input(({process_input[311:208]})), .process_output(inner2_0_process_output));
  dem #(.INSTANCE_NAME("inner3_0")) inner3_0(.CLK(CLK), .CE(process_CE), .process_input(({process_input[415:312]})), .process_output(inner3_0_process_output));
  dem #(.INSTANCE_NAME("inner4_0")) inner4_0(.CLK(CLK), .CE(process_CE), .process_input(({process_input[519:416]})), .process_output(inner4_0_process_output));
  dem #(.INSTANCE_NAME("inner5_0")) inner5_0(.CLK(CLK), .CE(process_CE), .process_input(({process_input[623:520]})), .process_output(inner5_0_process_output));
  dem #(.INSTANCE_NAME("inner6_0")) inner6_0(.CLK(CLK), .CE(process_CE), .process_input(({process_input[727:624]})), .process_output(inner6_0_process_output));
  dem #(.INSTANCE_NAME("inner7_0")) inner7_0(.CLK(CLK), .CE(process_CE), .process_input(({process_input[831:728]})), .process_output(inner7_0_process_output));
endmodule

module liftXYSeqPointwise_lambda(input CLK, input CE, input [831:0] process_input, output [191:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [831:0] unp_process_output;
  wire [191:0] f_process_output;
  assign process_output = f_process_output;
  // function: process pure=true delay=15
  // function: reset pure=true delay=0
  packTupleArrays_table__0x42bdcbb0 #(.INSTANCE_NAME("unp")) unp(.CLK(CLK), .process_CE(CE), .process_input(process_input), .process_output(unp_process_output));
  map_dem_W8_H1 #(.INSTANCE_NAME("f")) f(.CLK(CLK), .process_CE(CE), .process_input(unp_process_output), .process_output(f_process_output));
endmodule

module liftXYSeq_lambda(input CLK, input process_valid, input CE, input [575:0] process_input, output [191:0] process_output, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  wire [255:0] p_process_output;
  reg [575:0] process_input_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_input_delay1_validunnamednull0_CECE <= process_input; end end
  wire [191:0] m_process_output;
  assign process_output = m_process_output;
  // function: process pure=false delay=16
  // function: reset pure=false delay=0
  PosSeq_W656_H482_T8 #(.INSTANCE_NAME("p")) p(.CLK(CLK), .process_valid(process_valid), .CE(CE), .process_output(p_process_output), .reset(reset));
  liftXYSeqPointwise_lambda #(.INSTANCE_NAME("m")) m(.CLK(CLK), .CE(CE), .process_input({process_input_delay1_validunnamednull0_CECE,p_process_output}), .process_output(m_process_output));
endmodule

module demtop(input CLK, input process_valid, input CE, input [63:0] process_input, output [191:0] process_output, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  wire [239:0] st_process_output;
  wire [575:0] convstencils_process_output;
  reg process_valid_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay1_validunnamednull0_CECE <= process_valid; end end
  reg process_valid_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay2_validunnamednull0_CECE <= process_valid_delay1_validunnamednull0_CECE; end end
  wire [191:0] dem_process_output;
  assign process_output = dem_process_output;
  // function: process pure=false delay=18
  // function: reset pure=false delay=0
  stencilLinebuffer_Auint8_w656_h482_xmin2_ymin2 #(.INSTANCE_NAME("st")) st(.CLK(CLK), .process_valid(process_valid), .CE(CE), .process_input(process_input), .process_output(st_process_output), .reset(reset));
  unpackStencil_W3_H3_T8 #(.INSTANCE_NAME("convstencils")) convstencils(.CLK(CLK), .process_CE(CE), .inp(st_process_output), .process_output(convstencils_process_output));
  liftXYSeq_lambda #(.INSTANCE_NAME("dem")) dem(.CLK(CLK), .process_valid(process_valid_delay2_validunnamednull0_CECE), .CE(CE), .process_input(convstencils_process_output), .process_output(dem_process_output), .reset(reset));
endmodule

module ccm(input CLK, input process_CE, input [23:0] ccminp, output [23:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] unnamedcast4947USEDMULTIPLEcast = {8'b0,(8'd185)};
  wire [15:0] unnamedcast4948USEDMULTIPLEcast = {8'b0,({ccminp[7:0]})};
  reg [15:0] unnamedbinop4949_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop4949_delay1_validunnamednull0_CEprocess_CE <= {(unnamedcast4947USEDMULTIPLEcast*unnamedcast4948USEDMULTIPLEcast)}; end end
  wire [15:0] unnamedcast4953USEDMULTIPLEcast = {8'b0,(8'd0)};
  wire [15:0] unnamedcast4954USEDMULTIPLEcast = {8'b0,({ccminp[15:8]})};
  reg [15:0] unnamedbinop4955_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop4955_delay1_validunnamednull0_CEprocess_CE <= {(unnamedcast4953USEDMULTIPLEcast*unnamedcast4954USEDMULTIPLEcast)}; end end
  wire [16:0] unnamedcast4957USEDMULTIPLEcast = {1'b0,unnamedbinop4955_delay1_validunnamednull0_CEprocess_CE};
  reg [16:0] unnamedbinop4958_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop4958_delay1_validunnamednull0_CEprocess_CE <= {({1'b0,unnamedbinop4949_delay1_validunnamednull0_CEprocess_CE}+unnamedcast4957USEDMULTIPLEcast)}; end end
  wire [15:0] unnamedcast4963USEDMULTIPLEcast = {8'b0,({ccminp[23:16]})};
  reg [15:0] unnamedbinop4964_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop4964_delay1_validunnamednull0_CEprocess_CE <= {(unnamedcast4953USEDMULTIPLEcast*unnamedcast4963USEDMULTIPLEcast)}; end end
  reg [17:0] unnamedcast4966_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast4966_delay1_validunnamednull0_CEprocess_CE <= {2'b0,unnamedbinop4964_delay1_validunnamednull0_CEprocess_CE}; end end
  reg [17:0] unnamedbinop4967_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop4967_delay1_validunnamednull0_CEprocess_CE <= {({1'b0,unnamedbinop4958_delay1_validunnamednull0_CEprocess_CE}+unnamedcast4966_delay1_validunnamednull0_CEprocess_CE)}; end end
  reg [17:0] unnamedcast4969_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast4969_delay1_validunnamednull0_CEprocess_CE <= (18'd7); end end
  reg [17:0] unnamedcast4969_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast4969_delay2_validunnamednull0_CEprocess_CE <= unnamedcast4969_delay1_validunnamednull0_CEprocess_CE; end end
  reg [17:0] unnamedcast4969_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast4969_delay3_validunnamednull0_CEprocess_CE <= unnamedcast4969_delay2_validunnamednull0_CEprocess_CE; end end
  reg [17:0] unnamedbinop4970_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop4970_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop4967_delay1_validunnamednull0_CEprocess_CE>>>unnamedcast4969_delay3_validunnamednull0_CEprocess_CE)}; end end
  wire [10:0] unnamedcast4971USEDMULTIPLEcast = unnamedbinop4970_delay1_validunnamednull0_CEprocess_CE[10:0];
  reg [10:0] unnamedcast4973_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast4973_delay1_validunnamednull0_CEprocess_CE <= {3'b0,(8'd255)}; end end
  reg [10:0] unnamedcast4973_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast4973_delay2_validunnamednull0_CEprocess_CE <= unnamedcast4973_delay1_validunnamednull0_CEprocess_CE; end end
  reg [10:0] unnamedcast4973_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast4973_delay3_validunnamednull0_CEprocess_CE <= unnamedcast4973_delay2_validunnamednull0_CEprocess_CE; end end
  reg [10:0] unnamedcast4973_delay4_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast4973_delay4_validunnamednull0_CEprocess_CE <= unnamedcast4973_delay3_validunnamednull0_CEprocess_CE; end end
  reg unnamedbinop4974_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop4974_delay1_validunnamednull0_CEprocess_CE <= {((unnamedcast4971USEDMULTIPLEcast)>(unnamedcast4973_delay4_validunnamednull0_CEprocess_CE))}; end end
  reg [10:0] unnamedcast4976_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast4976_delay1_validunnamednull0_CEprocess_CE <= (11'd255); end end
  reg [10:0] unnamedcast4976_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast4976_delay2_validunnamednull0_CEprocess_CE <= unnamedcast4976_delay1_validunnamednull0_CEprocess_CE; end end
  reg [10:0] unnamedcast4976_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast4976_delay3_validunnamednull0_CEprocess_CE <= unnamedcast4976_delay2_validunnamednull0_CEprocess_CE; end end
  reg [10:0] unnamedcast4976_delay4_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast4976_delay4_validunnamednull0_CEprocess_CE <= unnamedcast4976_delay3_validunnamednull0_CEprocess_CE; end end
  reg [10:0] unnamedcast4976_delay5_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast4976_delay5_validunnamednull0_CEprocess_CE <= unnamedcast4976_delay4_validunnamednull0_CEprocess_CE; end end
  reg [10:0] unnamedcast4971_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast4971_delay1_validunnamednull0_CEprocess_CE <= unnamedcast4971USEDMULTIPLEcast; end end
  reg [10:0] unnamedselect4977_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedselect4977_delay1_validunnamednull0_CEprocess_CE <= ((unnamedbinop4974_delay1_validunnamednull0_CEprocess_CE)?(unnamedcast4976_delay5_validunnamednull0_CEprocess_CE):(unnamedcast4971_delay1_validunnamednull0_CEprocess_CE)); end end
  reg [15:0] unnamedbinop4984_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop4984_delay1_validunnamednull0_CEprocess_CE <= {(unnamedcast4953USEDMULTIPLEcast*unnamedcast4948USEDMULTIPLEcast)}; end end
  wire [16:0] unnamedcast4991USEDMULTIPLEcast = {1'b0,unnamedbinop4984_delay1_validunnamednull0_CEprocess_CE};
  reg [15:0] unnamedbinop4990_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop4990_delay1_validunnamednull0_CEprocess_CE <= {({8'b0,(8'd145)}*unnamedcast4954USEDMULTIPLEcast)}; end end
  reg [16:0] unnamedbinop4993_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop4993_delay1_validunnamednull0_CEprocess_CE <= {(unnamedcast4991USEDMULTIPLEcast+{1'b0,unnamedbinop4990_delay1_validunnamednull0_CEprocess_CE})}; end end
  reg [17:0] unnamedbinop5002_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop5002_delay1_validunnamednull0_CEprocess_CE <= {({1'b0,unnamedbinop4993_delay1_validunnamednull0_CEprocess_CE}+unnamedcast4966_delay1_validunnamednull0_CEprocess_CE)}; end end
  reg [17:0] unnamedbinop5005_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop5005_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop5002_delay1_validunnamednull0_CEprocess_CE>>>unnamedcast4969_delay3_validunnamednull0_CEprocess_CE)}; end end
  wire [10:0] unnamedcast5006USEDMULTIPLEcast = unnamedbinop5005_delay1_validunnamednull0_CEprocess_CE[10:0];
  reg unnamedbinop5009_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop5009_delay1_validunnamednull0_CEprocess_CE <= {((unnamedcast5006USEDMULTIPLEcast)>(unnamedcast4973_delay4_validunnamednull0_CEprocess_CE))}; end end
  reg [10:0] unnamedcast5006_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast5006_delay1_validunnamednull0_CEprocess_CE <= unnamedcast5006USEDMULTIPLEcast; end end
  reg [10:0] unnamedselect5012_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedselect5012_delay1_validunnamednull0_CEprocess_CE <= ((unnamedbinop5009_delay1_validunnamednull0_CEprocess_CE)?(unnamedcast4976_delay5_validunnamednull0_CEprocess_CE):(unnamedcast5006_delay1_validunnamednull0_CEprocess_CE)); end end
  reg [16:0] unnamedbinop5028_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop5028_delay1_validunnamednull0_CEprocess_CE <= {(unnamedcast4991USEDMULTIPLEcast+unnamedcast4957USEDMULTIPLEcast)}; end end
  reg [15:0] unnamedbinop5034_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop5034_delay1_validunnamednull0_CEprocess_CE <= {(unnamedcast4947USEDMULTIPLEcast*unnamedcast4963USEDMULTIPLEcast)}; end end
  reg [17:0] unnamedcast5036_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast5036_delay1_validunnamednull0_CEprocess_CE <= {2'b0,unnamedbinop5034_delay1_validunnamednull0_CEprocess_CE}; end end
  reg [17:0] unnamedbinop5037_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop5037_delay1_validunnamednull0_CEprocess_CE <= {({1'b0,unnamedbinop5028_delay1_validunnamednull0_CEprocess_CE}+unnamedcast5036_delay1_validunnamednull0_CEprocess_CE)}; end end
  reg [17:0] unnamedbinop5040_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop5040_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop5037_delay1_validunnamednull0_CEprocess_CE>>>unnamedcast4969_delay3_validunnamednull0_CEprocess_CE)}; end end
  wire [10:0] unnamedcast5041USEDMULTIPLEcast = unnamedbinop5040_delay1_validunnamednull0_CEprocess_CE[10:0];
  reg unnamedbinop5044_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop5044_delay1_validunnamednull0_CEprocess_CE <= {((unnamedcast5041USEDMULTIPLEcast)>(unnamedcast4973_delay4_validunnamednull0_CEprocess_CE))}; end end
  reg [10:0] unnamedcast5041_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast5041_delay1_validunnamednull0_CEprocess_CE <= unnamedcast5041USEDMULTIPLEcast; end end
  reg [10:0] unnamedselect5047_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedselect5047_delay1_validunnamednull0_CEprocess_CE <= ((unnamedbinop5044_delay1_validunnamednull0_CEprocess_CE)?(unnamedcast4976_delay5_validunnamednull0_CEprocess_CE):(unnamedcast5041_delay1_validunnamednull0_CEprocess_CE)); end end
  assign process_output = {unnamedselect5047_delay1_validunnamednull0_CEprocess_CE[7:0],unnamedselect5012_delay1_validunnamednull0_CEprocess_CE[7:0],unnamedselect4977_delay1_validunnamednull0_CEprocess_CE[7:0]};
  // function: process pure=true delay=6
endmodule

module map_ccm_W8_H1(input CLK, input process_CE, input [191:0] process_input, output [191:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [23:0] inner0_0_process_output;
  wire [23:0] inner1_0_process_output;
  wire [23:0] inner2_0_process_output;
  wire [23:0] inner3_0_process_output;
  wire [23:0] inner4_0_process_output;
  wire [23:0] inner5_0_process_output;
  wire [23:0] inner6_0_process_output;
  wire [23:0] inner7_0_process_output;
  assign process_output = {inner7_0_process_output,inner6_0_process_output,inner5_0_process_output,inner4_0_process_output,inner3_0_process_output,inner2_0_process_output,inner1_0_process_output,inner0_0_process_output};
  // function: process pure=true delay=6
  ccm #(.INSTANCE_NAME("inner0_0")) inner0_0(.CLK(CLK), .process_CE(process_CE), .ccminp(({process_input[23:0]})), .process_output(inner0_0_process_output));
  ccm #(.INSTANCE_NAME("inner1_0")) inner1_0(.CLK(CLK), .process_CE(process_CE), .ccminp(({process_input[47:24]})), .process_output(inner1_0_process_output));
  ccm #(.INSTANCE_NAME("inner2_0")) inner2_0(.CLK(CLK), .process_CE(process_CE), .ccminp(({process_input[71:48]})), .process_output(inner2_0_process_output));
  ccm #(.INSTANCE_NAME("inner3_0")) inner3_0(.CLK(CLK), .process_CE(process_CE), .ccminp(({process_input[95:72]})), .process_output(inner3_0_process_output));
  ccm #(.INSTANCE_NAME("inner4_0")) inner4_0(.CLK(CLK), .process_CE(process_CE), .ccminp(({process_input[119:96]})), .process_output(inner4_0_process_output));
  ccm #(.INSTANCE_NAME("inner5_0")) inner5_0(.CLK(CLK), .process_CE(process_CE), .ccminp(({process_input[143:120]})), .process_output(inner5_0_process_output));
  ccm #(.INSTANCE_NAME("inner6_0")) inner6_0(.CLK(CLK), .process_CE(process_CE), .ccminp(({process_input[167:144]})), .process_output(inner6_0_process_output));
  ccm #(.INSTANCE_NAME("inner7_0")) inner7_0(.CLK(CLK), .process_CE(process_CE), .ccminp(({process_input[191:168]})), .process_output(inner7_0_process_output));
endmodule

module bramSDP_WAROtrue_size256_bw1_obw1_CEtrue_inittable__0x403e5208(input CLK, input [7:0] inpRead, output [7:0] READ_OUT, input writeAndReturnOriginal_valid, input writeAndReturnOriginal_CE, input [15:0] inp, output [7:0] WARO_OUT);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(writeAndReturnOriginal_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'writeAndReturnOriginal'", INSTANCE_NAME);  end end
  wire [10:0] unnamedcast5244USEDMULTIPLEcast = {3'b0,(inp[7:0])};
  wire [7:0] bram_0_READ_OUTPUT;
  assign READ_OUT = {bram_0_READ_OUTPUT};
  wire [7:0] unnamedcast5239 = (inp[15:8]); // wire for bitslice
  wire [7:0] bram_0_SET_AND_RETURN_ORIG_OUTPUT;
  assign WARO_OUT = {bram_0_SET_AND_RETURN_ORIG_OUTPUT};
  // function: read pure=true delay=1
  // function: writeAndReturnOriginal pure=false delay=1
  reg [7:0] bram_0_DI_B;
reg [10:0] bram_0_addr_B;
wire [7:0] bram_0_DO_B;
wire [18:0] bram_0_INPUT;
assign bram_0_INPUT = {unnamedcast5239[7:0],unnamedcast5244USEDMULTIPLEcast};
RAMB16_S9_S9 #(.WRITE_MODE_A("READ_FIRST"),.WRITE_MODE_B("READ_FIRST"),.INIT_00(256'h2c2a29282726242322211f1e1d1b1a191816151312110f0e0c0b090706040200),.INIT_01(256'h4f4e4d4c4b4a4948474544434241403f3e3d3c3a3938373635343331302f2e2d),.INIT_02(256'h6f6f6e6d6c6b6a696867666564636261605f5e5c5b5a59585756555453525150),.INIT_03(256'h8e8d8c8b8a89898887868584838281807f7e7d7c7b7a79787776757473727170),.INIT_04(256'hacabaaa9a8a7a6a5a4a3a2a2a1a09f9e9d9c9b9a99989797969594939291908f),.INIT_05(256'hc8c7c6c5c4c4c3c2c1c0bfbebdbcbcbbbab9b8b7b6b5b4b4b3b2b1b0afaeadac),.INIT_06(256'he4e3e2e1e0dfdededddcdbdad9d8d8d7d6d5d4d3d2d1d1d0cfcecdcccbcbcac9),.INIT_07(256'hfffefdfcfbfaf9f9f8f7f6f5f4f4f3f2f1f0efefeeedecebeae9e9e8e7e6e5e4),.INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)) bram_0 (
.DIPA(1'b0),
.DIPB(1'b0),
.DIA(bram_0_INPUT[18:11]),
.DIB(bram_0_DI_B),
.DOA(bram_0_SET_AND_RETURN_ORIG_OUTPUT),
.DOB(bram_0_READ_OUTPUT),
.ADDRA(bram_0_INPUT[10:0]),
.ADDRB(unnamedcast5244USEDMULTIPLEcast),
.WEA(writeAndReturnOriginal_valid),
.WEB(1'd0),
.ENA(writeAndReturnOriginal_CE),
.ENB(writeAndReturnOriginal_CE),
.CLKA(CLK),
.CLKB(CLK),
.SSRA(1'b0),
.SSRB(1'b0)
);


endmodule

module LUT(input CLK, input process_valid, input process_CE, input [7:0] process_input, output [7:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  wire [7:0] LUT_READ_OUT;
  wire [7:0] LUT_WARO_OUT;
  assign process_output = LUT_READ_OUT;
  // function: process pure=false delay=1
  bramSDP_WAROtrue_size256_bw1_obw1_CEtrue_inittable__0x403e5208 #(.INSTANCE_NAME("LUT")) LUT(.CLK(CLK), .inpRead(process_input), .READ_OUT(LUT_READ_OUT), .writeAndReturnOriginal_valid({((1'd0)&&process_valid)}), .writeAndReturnOriginal_CE(process_CE), .inp({(8'd0),process_input}), .WARO_OUT(LUT_WARO_OUT));
endmodule

module map_LUT_W3_H1(input CLK, input process_valid, input process_CE, input [23:0] process_input, output [23:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  wire [7:0] inner0_0_process_output;
  wire [7:0] inner1_0_process_output;
  wire [7:0] inner2_0_process_output;
  assign process_output = {inner2_0_process_output,inner1_0_process_output,inner0_0_process_output};
  // function: process pure=false delay=1
  LUT #(.INSTANCE_NAME("inner0_0")) inner0_0(.CLK(CLK), .process_valid(process_valid), .process_CE(process_CE), .process_input(({process_input[7:0]})), .process_output(inner0_0_process_output));
  LUT #(.INSTANCE_NAME("inner1_0")) inner1_0(.CLK(CLK), .process_valid(process_valid), .process_CE(process_CE), .process_input(({process_input[15:8]})), .process_output(inner1_0_process_output));
  LUT #(.INSTANCE_NAME("inner2_0")) inner2_0(.CLK(CLK), .process_valid(process_valid), .process_CE(process_CE), .process_input(({process_input[23:16]})), .process_output(inner2_0_process_output));
endmodule

module map_map_LUT_W3_H1_W8_H1(input CLK, input process_valid, input process_CE, input [191:0] process_input, output [191:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  wire [23:0] inner0_0_process_output;
  wire [23:0] inner1_0_process_output;
  wire [23:0] inner2_0_process_output;
  wire [23:0] inner3_0_process_output;
  wire [23:0] inner4_0_process_output;
  wire [23:0] inner5_0_process_output;
  wire [23:0] inner6_0_process_output;
  wire [23:0] inner7_0_process_output;
  assign process_output = {inner7_0_process_output,inner6_0_process_output,inner5_0_process_output,inner4_0_process_output,inner3_0_process_output,inner2_0_process_output,inner1_0_process_output,inner0_0_process_output};
  // function: process pure=false delay=1
  map_LUT_W3_H1 #(.INSTANCE_NAME("inner0_0")) inner0_0(.CLK(CLK), .process_valid(process_valid), .process_CE(process_CE), .process_input(({process_input[23:0]})), .process_output(inner0_0_process_output));
  map_LUT_W3_H1 #(.INSTANCE_NAME("inner1_0")) inner1_0(.CLK(CLK), .process_valid(process_valid), .process_CE(process_CE), .process_input(({process_input[47:24]})), .process_output(inner1_0_process_output));
  map_LUT_W3_H1 #(.INSTANCE_NAME("inner2_0")) inner2_0(.CLK(CLK), .process_valid(process_valid), .process_CE(process_CE), .process_input(({process_input[71:48]})), .process_output(inner2_0_process_output));
  map_LUT_W3_H1 #(.INSTANCE_NAME("inner3_0")) inner3_0(.CLK(CLK), .process_valid(process_valid), .process_CE(process_CE), .process_input(({process_input[95:72]})), .process_output(inner3_0_process_output));
  map_LUT_W3_H1 #(.INSTANCE_NAME("inner4_0")) inner4_0(.CLK(CLK), .process_valid(process_valid), .process_CE(process_CE), .process_input(({process_input[119:96]})), .process_output(inner4_0_process_output));
  map_LUT_W3_H1 #(.INSTANCE_NAME("inner5_0")) inner5_0(.CLK(CLK), .process_valid(process_valid), .process_CE(process_CE), .process_input(({process_input[143:120]})), .process_output(inner5_0_process_output));
  map_LUT_W3_H1 #(.INSTANCE_NAME("inner6_0")) inner6_0(.CLK(CLK), .process_valid(process_valid), .process_CE(process_CE), .process_input(({process_input[167:144]})), .process_output(inner6_0_process_output));
  map_LUT_W3_H1 #(.INSTANCE_NAME("inner7_0")) inner7_0(.CLK(CLK), .process_valid(process_valid), .process_CE(process_CE), .process_input(({process_input[191:168]})), .process_output(inner7_0_process_output));
endmodule

module addChan(input CLK, input process_CE, input [23:0] inp, output [31:0] process_output);
parameter INSTANCE_NAME="INST";
  assign process_output = {(8'd0),({inp[23:16]}),({inp[15:8]}),({inp[7:0]})};
  // function: process pure=true delay=0
endmodule

module map_addChan_W8_H1(input CLK, input process_CE, input [191:0] process_input, output [255:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [31:0] inner0_0_process_output;
  wire [31:0] inner1_0_process_output;
  wire [31:0] inner2_0_process_output;
  wire [31:0] inner3_0_process_output;
  wire [31:0] inner4_0_process_output;
  wire [31:0] inner5_0_process_output;
  wire [31:0] inner6_0_process_output;
  wire [31:0] inner7_0_process_output;
  assign process_output = {inner7_0_process_output,inner6_0_process_output,inner5_0_process_output,inner4_0_process_output,inner3_0_process_output,inner2_0_process_output,inner1_0_process_output,inner0_0_process_output};
  // function: process pure=true delay=0
  addChan #(.INSTANCE_NAME("inner0_0")) inner0_0(.CLK(CLK), .process_CE(process_CE), .inp(({process_input[23:0]})), .process_output(inner0_0_process_output));
  addChan #(.INSTANCE_NAME("inner1_0")) inner1_0(.CLK(CLK), .process_CE(process_CE), .inp(({process_input[47:24]})), .process_output(inner1_0_process_output));
  addChan #(.INSTANCE_NAME("inner2_0")) inner2_0(.CLK(CLK), .process_CE(process_CE), .inp(({process_input[71:48]})), .process_output(inner2_0_process_output));
  addChan #(.INSTANCE_NAME("inner3_0")) inner3_0(.CLK(CLK), .process_CE(process_CE), .inp(({process_input[95:72]})), .process_output(inner3_0_process_output));
  addChan #(.INSTANCE_NAME("inner4_0")) inner4_0(.CLK(CLK), .process_CE(process_CE), .inp(({process_input[119:96]})), .process_output(inner4_0_process_output));
  addChan #(.INSTANCE_NAME("inner5_0")) inner5_0(.CLK(CLK), .process_CE(process_CE), .inp(({process_input[143:120]})), .process_output(inner5_0_process_output));
  addChan #(.INSTANCE_NAME("inner6_0")) inner6_0(.CLK(CLK), .process_CE(process_CE), .inp(({process_input[167:144]})), .process_output(inner6_0_process_output));
  addChan #(.INSTANCE_NAME("inner7_0")) inner7_0(.CLK(CLK), .process_CE(process_CE), .inp(({process_input[191:168]})), .process_output(inner7_0_process_output));
endmodule

module campipe(input CLK, input process_valid, input CE, input [63:0] process_input, output [255:0] process_output, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  wire [63:0] bl_process_output;
  reg process_valid_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay1_validunnamednull0_CECE <= process_valid; end end
  reg process_valid_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay2_validunnamednull0_CECE <= process_valid_delay1_validunnamednull0_CECE; end end
  reg process_valid_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay3_validunnamednull0_CECE <= process_valid_delay2_validunnamednull0_CECE; end end
  reg process_valid_delay4_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay4_validunnamednull0_CECE <= process_valid_delay3_validunnamednull0_CECE; end end
  reg process_valid_delay5_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay5_validunnamednull0_CECE <= process_valid_delay4_validunnamednull0_CECE; end end
  reg process_valid_delay6_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay6_validunnamednull0_CECE <= process_valid_delay5_validunnamednull0_CECE; end end
  wire [191:0] dem_process_output;
  wire [191:0] ccm_process_output;
  reg process_valid_delay7_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay7_validunnamednull0_CECE <= process_valid_delay6_validunnamednull0_CECE; end end
  reg process_valid_delay8_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay8_validunnamednull0_CECE <= process_valid_delay7_validunnamednull0_CECE; end end
  reg process_valid_delay9_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay9_validunnamednull0_CECE <= process_valid_delay8_validunnamednull0_CECE; end end
  reg process_valid_delay10_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay10_validunnamednull0_CECE <= process_valid_delay9_validunnamednull0_CECE; end end
  reg process_valid_delay11_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay11_validunnamednull0_CECE <= process_valid_delay10_validunnamednull0_CECE; end end
  reg process_valid_delay12_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay12_validunnamednull0_CECE <= process_valid_delay11_validunnamednull0_CECE; end end
  reg process_valid_delay13_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay13_validunnamednull0_CECE <= process_valid_delay12_validunnamednull0_CECE; end end
  reg process_valid_delay14_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay14_validunnamednull0_CECE <= process_valid_delay13_validunnamednull0_CECE; end end
  reg process_valid_delay15_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay15_validunnamednull0_CECE <= process_valid_delay14_validunnamednull0_CECE; end end
  reg process_valid_delay16_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay16_validunnamednull0_CECE <= process_valid_delay15_validunnamednull0_CECE; end end
  reg process_valid_delay17_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay17_validunnamednull0_CECE <= process_valid_delay16_validunnamednull0_CECE; end end
  reg process_valid_delay18_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay18_validunnamednull0_CECE <= process_valid_delay17_validunnamednull0_CECE; end end
  reg process_valid_delay19_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay19_validunnamednull0_CECE <= process_valid_delay18_validunnamednull0_CECE; end end
  reg process_valid_delay20_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay20_validunnamednull0_CECE <= process_valid_delay19_validunnamednull0_CECE; end end
  reg process_valid_delay21_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay21_validunnamednull0_CECE <= process_valid_delay20_validunnamednull0_CECE; end end
  reg process_valid_delay22_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay22_validunnamednull0_CECE <= process_valid_delay21_validunnamednull0_CECE; end end
  reg process_valid_delay23_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay23_validunnamednull0_CECE <= process_valid_delay22_validunnamednull0_CECE; end end
  reg process_valid_delay24_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay24_validunnamednull0_CECE <= process_valid_delay23_validunnamednull0_CECE; end end
  reg process_valid_delay25_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay25_validunnamednull0_CECE <= process_valid_delay24_validunnamednull0_CECE; end end
  reg process_valid_delay26_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay26_validunnamednull0_CECE <= process_valid_delay25_validunnamednull0_CECE; end end
  reg process_valid_delay27_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay27_validunnamednull0_CECE <= process_valid_delay26_validunnamednull0_CECE; end end
  reg process_valid_delay28_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay28_validunnamednull0_CECE <= process_valid_delay27_validunnamednull0_CECE; end end
  reg process_valid_delay29_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay29_validunnamednull0_CECE <= process_valid_delay28_validunnamednull0_CECE; end end
  reg process_valid_delay30_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay30_validunnamednull0_CECE <= process_valid_delay29_validunnamednull0_CECE; end end
  wire [191:0] gam_process_output;
  wire [255:0] addchan_process_output;
  assign process_output = addchan_process_output;
  // function: process pure=false delay=31
  // function: reset pure=false delay=0
  map_blackLevel_W8_H1 #(.INSTANCE_NAME("bl")) bl(.CLK(CLK), .process_CE(CE), .process_input(process_input), .process_output(bl_process_output));
  demtop #(.INSTANCE_NAME("dem")) dem(.CLK(CLK), .process_valid(process_valid_delay6_validunnamednull0_CECE), .CE(CE), .process_input(bl_process_output), .process_output(dem_process_output), .reset(reset));
  map_ccm_W8_H1 #(.INSTANCE_NAME("ccm")) ccm(.CLK(CLK), .process_CE(CE), .process_input(dem_process_output), .process_output(ccm_process_output));
  map_map_LUT_W3_H1_W8_H1 #(.INSTANCE_NAME("gam")) gam(.CLK(CLK), .process_valid(process_valid_delay30_validunnamednull0_CECE), .process_CE(CE), .process_input(ccm_process_output), .process_output(gam_process_output));
  map_addChan_W8_H1 #(.INSTANCE_NAME("addchan")) addchan(.CLK(CLK), .process_CE(CE), .process_input(gam_process_output), .process_output(addchan_process_output));
endmodule

module MakeHandshake_campipe(input CLK, input ready_downstream, output ready, input reset, input [64:0] process_input, output [256:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  assign ready = ready_downstream;
  wire unnamedbinop6208USEDMULTIPLEbinop = {(ready_downstream||reset)};
  wire unnamedcast6216USEDMULTIPLEcast = (process_input[64]);
  wire [255:0] inner_process_output;
  wire validBitDelay_campipe_pushPop_out;
  always @(posedge CLK) begin if({(~{(unnamedcast6216USEDMULTIPLEcast===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: MakeHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = {validBitDelay_campipe_pushPop_out,inner_process_output};
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  ShiftRegister_31_CEtrue_TY1 #(.INSTANCE_NAME("validBitDelay_campipe")) validBitDelay_campipe(.CLK(CLK), .pushPop_valid({(~reset)}), .CE(unnamedbinop6208USEDMULTIPLEbinop), .sr_input(unnamedcast6216USEDMULTIPLEcast), .pushPop_out(validBitDelay_campipe_pushPop_out), .reset(reset));
  campipe #(.INSTANCE_NAME("inner")) inner(.CLK(CLK), .process_valid(unnamedcast6216USEDMULTIPLEcast), .CE(unnamedbinop6208USEDMULTIPLEbinop), .process_input((process_input[63:0])), .process_output(inner_process_output), .reset(reset));
endmodule

module SSR_W8_H1_T8_Auint8_4_1_(input CLK, input process_valid, input process_CE, input [255:0] inp, output [479:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  reg [31:0] SR_x0_y0;
  reg [31:0] SR_x1_y0;
  reg [31:0] SR_x2_y0;
  reg [31:0] SR_x3_y0;
  reg [31:0] SR_x4_y0;
  reg [31:0] SR_x5_y0;
  reg [31:0] SR_x6_y0;
  wire [31:0] unnamedcast6234USEDMULTIPLEcast = ({inp[63:32]});
  wire [31:0] unnamedcast6232USEDMULTIPLEcast = ({inp[95:64]});
  wire [31:0] unnamedcast6230USEDMULTIPLEcast = ({inp[127:96]});
  wire [31:0] unnamedcast6228USEDMULTIPLEcast = ({inp[159:128]});
  wire [31:0] unnamedcast6226USEDMULTIPLEcast = ({inp[191:160]});
  wire [31:0] unnamedcast6224USEDMULTIPLEcast = ({inp[223:192]});
  wire [31:0] unnamedcast6222USEDMULTIPLEcast = ({inp[255:224]});
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x6_y0 <= unnamedcast6222USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x5_y0 <= unnamedcast6224USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x4_y0 <= unnamedcast6226USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x3_y0 <= unnamedcast6228USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x2_y0 <= unnamedcast6230USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x1_y0 <= unnamedcast6232USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x0_y0 <= unnamedcast6234USEDMULTIPLEcast; end end
  assign process_output = {unnamedcast6222USEDMULTIPLEcast,unnamedcast6224USEDMULTIPLEcast,unnamedcast6226USEDMULTIPLEcast,unnamedcast6228USEDMULTIPLEcast,unnamedcast6230USEDMULTIPLEcast,unnamedcast6232USEDMULTIPLEcast,unnamedcast6234USEDMULTIPLEcast,({inp[31:0]}),SR_x6_y0,SR_x5_y0,SR_x4_y0,SR_x3_y0,SR_x2_y0,SR_x1_y0,SR_x0_y0};
  // function: process pure=false delay=0
  // function: reset pure=true delay=0
endmodule

module slice_typeuint8_4_1__15_1__xl0_xh7_yl0_yh0(input CLK, input process_CE, input [479:0] inp, output [255:0] process_output);
parameter INSTANCE_NAME="INST";
  assign process_output = {({inp[255:224]}),({inp[223:192]}),({inp[191:160]}),({inp[159:128]}),({inp[127:96]}),({inp[95:64]}),({inp[63:32]}),({inp[31:0]})};
  // function: process pure=true delay=0
endmodule

module CropSeq_W656_H482_T8(input CLK, input process_CE, input [511:0] process_input, output [256:0] process_output);
parameter INSTANCE_NAME="INST";
  reg [255:0] unnamedcast6314_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast6314_delay1_validunnamednull0_CEprocess_CE <= (process_input[511:256]); end end
  reg [255:0] unnamedcast6314_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast6314_delay2_validunnamednull0_CEprocess_CE <= unnamedcast6314_delay1_validunnamednull0_CEprocess_CE; end end
  reg [255:0] unnamedcast6314_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast6314_delay3_validunnamednull0_CEprocess_CE <= unnamedcast6314_delay2_validunnamednull0_CEprocess_CE; end end
  wire [255:0] unnamedcast6316 = (process_input[255:0]); // wire for array index
  wire [31:0] unnamedcast6318USEDMULTIPLEcast = ({unnamedcast6316[31:0]});
  wire [15:0] unnamedcast6320USEDMULTIPLEcast = (unnamedcast6318USEDMULTIPLEcast[15:0]);
  reg unnamedbinop6332_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop6332_delay1_validunnamednull0_CEprocess_CE <= {((unnamedcast6320USEDMULTIPLEcast)>=((16'd16)))}; end end
  wire [15:0] unnamedcast6326USEDMULTIPLEcast = (unnamedcast6318USEDMULTIPLEcast[31:16]);
  reg unnamedbinop6334_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop6334_delay1_validunnamednull0_CEprocess_CE <= {((unnamedcast6326USEDMULTIPLEcast)>=((16'd2)))}; end end
  reg unnamedbinop6335_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop6335_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop6332_delay1_validunnamednull0_CEprocess_CE&&unnamedbinop6334_delay1_validunnamednull0_CEprocess_CE)}; end end
  reg unnamedbinop6337_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop6337_delay1_validunnamednull0_CEprocess_CE <= {((unnamedcast6320USEDMULTIPLEcast)<((16'd656)))}; end end
  reg unnamedbinop6339_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop6339_delay1_validunnamednull0_CEprocess_CE <= {((unnamedcast6326USEDMULTIPLEcast)<((16'd482)))}; end end
  reg unnamedbinop6340_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop6340_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop6337_delay1_validunnamednull0_CEprocess_CE&&unnamedbinop6339_delay1_validunnamednull0_CEprocess_CE)}; end end
  reg unnamedbinop6341_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop6341_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop6335_delay1_validunnamednull0_CEprocess_CE&&unnamedbinop6340_delay1_validunnamednull0_CEprocess_CE)}; end end
  assign process_output = {unnamedbinop6341_delay1_validunnamednull0_CEprocess_CE,unnamedcast6314_delay3_validunnamednull0_CEprocess_CE};
  // function: process pure=true delay=3
endmodule

module liftXYSeq_lift_CropSeq_W656_H482_T8(input CLK, input process_valid, input CE, input [255:0] process_input, output [256:0] process_output, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  wire [255:0] p_process_output;
  reg [255:0] process_input_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_input_delay1_validunnamednull0_CECE <= process_input; end end
  wire [256:0] m_process_output;
  assign process_output = m_process_output;
  // function: process pure=false delay=4
  // function: reset pure=false delay=0
  PosSeq_W656_H482_T8 #(.INSTANCE_NAME("p")) p(.CLK(CLK), .process_valid(process_valid), .CE(CE), .process_output(p_process_output), .reset(reset));
  CropSeq_W656_H482_T8 #(.INSTANCE_NAME("m")) m(.CLK(CLK), .process_CE(CE), .process_input({process_input_delay1_validunnamednull0_CECE,p_process_output}), .process_output(m_process_output));
endmodule

module cropHelperSeq(input CLK, input process_valid, input CE, input [255:0] process_input, output [256:0] process_output, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  wire [479:0] SSR_process_output;
  wire [255:0] slice_process_output;
  wire [256:0] crop_process_output;
  assign process_output = crop_process_output;
  // function: process pure=false delay=4
  // function: reset pure=false delay=0
  SSR_W8_H1_T8_Auint8_4_1_ #(.INSTANCE_NAME("SSR")) SSR(.CLK(CLK), .process_valid(process_valid), .process_CE(CE), .inp(process_input), .process_output(SSR_process_output));
  slice_typeuint8_4_1__15_1__xl0_xh7_yl0_yh0 #(.INSTANCE_NAME("slice")) slice(.CLK(CLK), .process_CE(CE), .inp(SSR_process_output), .process_output(slice_process_output));
  liftXYSeq_lift_CropSeq_W656_H482_T8 #(.INSTANCE_NAME("crop")) crop(.CLK(CLK), .process_valid(process_valid), .CE(CE), .process_input(slice_process_output), .process_output(crop_process_output), .reset(reset));
endmodule

module LiftDecimate_cropHelperSeq(input CLK, output ready, input reset, input CE, input process_valid, input [256:0] process_input, output [256:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  assign ready = (1'd1);
  wire unnamedcast6515USEDMULTIPLEcast = (process_input[256]);
  wire [256:0] LiftDecimate_inner_cropHelperSeq_process_output;
  reg [255:0] unnamedcast6518_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast6518_delay1_validunnamednull0_CECE <= (LiftDecimate_inner_cropHelperSeq_process_output[255:0]); end end
  reg unnamedcast6515_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast6515_delay1_validunnamednull0_CECE <= unnamedcast6515USEDMULTIPLEcast; end end
  reg unnamedcast6515_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast6515_delay2_validunnamednull0_CECE <= unnamedcast6515_delay1_validunnamednull0_CECE; end end
  reg unnamedcast6515_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast6515_delay3_validunnamednull0_CECE <= unnamedcast6515_delay2_validunnamednull0_CECE; end end
  reg unnamedcast6515_delay4_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast6515_delay4_validunnamednull0_CECE <= unnamedcast6515_delay3_validunnamednull0_CECE; end end
  reg unnamedbinop6523_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedbinop6523_delay1_validunnamednull0_CECE <= {((LiftDecimate_inner_cropHelperSeq_process_output[256])&&unnamedcast6515_delay4_validunnamednull0_CECE)}; end end
  assign process_output = {unnamedbinop6523_delay1_validunnamednull0_CECE,unnamedcast6518_delay1_validunnamednull0_CECE};
  // function: ready pure=true delay=0
  // function: reset pure=false delay=0
  // function: process pure=false delay=5
  cropHelperSeq #(.INSTANCE_NAME("LiftDecimate_inner_cropHelperSeq")) LiftDecimate_inner_cropHelperSeq(.CLK(CLK), .process_valid({(unnamedcast6515USEDMULTIPLEcast&&process_valid)}), .CE(CE), .process_input((process_input[255:0])), .process_output(LiftDecimate_inner_cropHelperSeq_process_output), .reset(reset));
endmodule

module ShiftRegister_5_CEtrue_TY1(input CLK, input pushPop_valid, input CE, input sr_input, output pushPop_out, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'pushPop'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  reg SR5;
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR1' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR1' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR1' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6626USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(sr_input):((1'd0)))};
  reg SR1;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6626USEDMULTIPLEcallArbitrate[1]) && CE) begin SR1 <= (unnamedcallArbitrate6626USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR2' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR2' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR2' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6632USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR1):((1'd0)))};
  reg SR2;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6632USEDMULTIPLEcallArbitrate[1]) && CE) begin SR2 <= (unnamedcallArbitrate6632USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR3' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR3' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR3' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6638USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR2):((1'd0)))};
  reg SR3;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6638USEDMULTIPLEcallArbitrate[1]) && CE) begin SR3 <= (unnamedcallArbitrate6638USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR4' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR4' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR4' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6644USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR3):((1'd0)))};
  reg SR4;  always @ (posedge CLK) begin if ((unnamedcallArbitrate6644USEDMULTIPLEcallArbitrate[1]) && CE) begin SR4 <= (unnamedcallArbitrate6644USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR5' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR5' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR5' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate6650USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR4):((1'd0)))};
    always @ (posedge CLK) begin if ((unnamedcallArbitrate6650USEDMULTIPLEcallArbitrate[1]) && CE) begin SR5 <= (unnamedcallArbitrate6650USEDMULTIPLEcallArbitrate[0]); end end
  assign pushPop_out = SR5;
  // function: pushPop pure=false delay=0
  // function: reset pure=false delay=0
endmodule

module LiftHandshake_LiftDecimate_cropHelperSeq(input CLK, input ready_downstream, output ready, input reset, input [256:0] process_input, output [256:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire inner_LiftDecimate_cropHelperSeq_ready;
  assign ready = {(inner_LiftDecimate_cropHelperSeq_ready&&ready_downstream)};
  wire unnamedbinop6563USEDMULTIPLEbinop = {(reset||ready_downstream)};
  wire unnamedunary6564USEDMULTIPLEunary = {(~reset)};
  wire [256:0] inner_LiftDecimate_cropHelperSeq_process_output;
  wire validBitDelay_LiftDecimate_cropHelperSeq_pushPop_out;
  wire [256:0] unnamedtuple6664USEDMULTIPLEtuple = {{((inner_LiftDecimate_cropHelperSeq_process_output[256])&&validBitDelay_LiftDecimate_cropHelperSeq_pushPop_out)},(inner_LiftDecimate_cropHelperSeq_process_output[255:0])};
  always @(posedge CLK) begin if({(~{((unnamedtuple6664USEDMULTIPLEtuple[256])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: output valid bit should not be X!",INSTANCE_NAME); end end
  always @(posedge CLK) begin if({(~{((process_input[256])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = unnamedtuple6664USEDMULTIPLEtuple;
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  LiftDecimate_cropHelperSeq #(.INSTANCE_NAME("inner_LiftDecimate_cropHelperSeq")) inner_LiftDecimate_cropHelperSeq(.CLK(CLK), .ready(inner_LiftDecimate_cropHelperSeq_ready), .reset(reset), .CE(unnamedbinop6563USEDMULTIPLEbinop), .process_valid(unnamedunary6564USEDMULTIPLEunary), .process_input(process_input), .process_output(inner_LiftDecimate_cropHelperSeq_process_output));
  ShiftRegister_5_CEtrue_TY1 #(.INSTANCE_NAME("validBitDelay_LiftDecimate_cropHelperSeq")) validBitDelay_LiftDecimate_cropHelperSeq(.CLK(CLK), .pushPop_valid(unnamedunary6564USEDMULTIPLEunary), .CE(unnamedbinop6563USEDMULTIPLEbinop), .sr_input((1'd1)), .pushPop_out(validBitDelay_LiftDecimate_cropHelperSeq_pushPop_out), .reset(reset));
endmodule

module hsfn(input CLK, input ready_downstream, output ready, input reset, input [64:0] process_input, output [256:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire [2:0] unnamedtuple12189USEDMULTIPLEtuple = {(1'd1),(1'd1),ready_downstream};
  wire f1_store_ready;
  wire pad_ready;
  wire f2_store_ready;
  wire crop_ready;
  wire HH_ready;
  wire f1_load_ready;
  wire f2_load_ready;
  assign ready = pad_ready;
  wire [0:0] unnamedtuple12159USEDMULTIPLEtuple = {(1'd1)};
  wire [256:0] f2_load_output;
  wire [64:0] pad_process_output;
  wire [0:0] f1_store_output;
  wire [64:0] f1_load_output;
  wire [256:0] HH_process_output;
  wire [256:0] crop_process_output;
  wire [0:0] f2_store_output;
  assign process_output = f2_load_output;
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  LiftHandshake_RunIffReady_LiftDecimate_fifo_128_uint8_8_1_ #(.INSTANCE_NAME("f1")) f1(.CLK(CLK), .load_input(unnamedtuple12159USEDMULTIPLEtuple), .load_output(f1_load_output), .store_reset(reset), .store_ready_downstream((unnamedtuple12189USEDMULTIPLEtuple[1])), .store_ready(f1_store_ready), .load_ready_downstream(HH_ready), .load_ready(f1_load_ready), .load_reset(reset), .store_input(pad_process_output), .store_output(f1_store_output));
  LiftHandshake_RunIffReady_LiftDecimate_fifo_128_uint8_4_1__8_1_ #(.INSTANCE_NAME("f2")) f2(.CLK(CLK), .load_input(unnamedtuple12159USEDMULTIPLEtuple), .load_output(f2_load_output), .store_reset(reset), .store_ready_downstream((unnamedtuple12189USEDMULTIPLEtuple[2])), .store_ready(f2_store_ready), .load_ready_downstream((unnamedtuple12189USEDMULTIPLEtuple[0])), .load_ready(f2_load_ready), .load_reset(reset), .store_input(crop_process_output), .store_output(f2_store_output));
  LiftHandshake_WaitOnInput_PadSeq_W640_H480_L8_R8_B1_Top1_T88 #(.INSTANCE_NAME("pad")) pad(.CLK(CLK), .ready_downstream(f1_store_ready), .ready(pad_ready), .reset(reset), .process_input(process_input), .process_output(pad_process_output));
  MakeHandshake_campipe #(.INSTANCE_NAME("HH")) HH(.CLK(CLK), .ready_downstream(crop_ready), .ready(HH_ready), .reset(reset), .process_input(f1_load_output), .process_output(HH_process_output));
  LiftHandshake_LiftDecimate_cropHelperSeq #(.INSTANCE_NAME("crop")) crop(.CLK(CLK), .ready_downstream(f2_store_ready), .ready(crop_ready), .reset(reset), .process_input(HH_process_output), .process_output(crop_process_output));
endmodule

module sumwrap_uint16_to3(input CLK, input CE, input [31:0] process_input, output [15:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] unnamedcast12212USEDMULTIPLEcast = (process_input[15:0]);
  assign process_output = (({(unnamedcast12212USEDMULTIPLEcast==(16'd3))})?((16'd0)):({(unnamedcast12212USEDMULTIPLEcast+(process_input[31:16]))}));
  // function: process pure=true delay=0
endmodule

module RegBy_sumwrap_uint16_to3_CEtrue_initnil(input CLK, input set_valid, input CE, input [15:0] set_inp, input setby_valid, input [15:0] setby_inp, output [15:0] SETBY_OUTPUT, output [15:0] GET_OUTPUT);
parameter INSTANCE_NAME="INST";
  reg [15:0] R;
  wire [15:0] regby_inner_process_output;
  always @(posedge CLK) begin if(set_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(setby_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,set_valid})+({4'b0,setby_valid})) > 5'd1) begin $display("error, function 'set' on instance 'R' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [16:0] unnamedcallArbitrate12252USEDMULTIPLEcallArbitrate = {(set_valid||setby_valid),((set_valid)?(set_inp):(regby_inner_process_output))};
    always @ (posedge CLK) begin if ((unnamedcallArbitrate12252USEDMULTIPLEcallArbitrate[16]) && CE) begin R <= (unnamedcallArbitrate12252USEDMULTIPLEcallArbitrate[15:0]); end end
  assign SETBY_OUTPUT = regby_inner_process_output;
  assign GET_OUTPUT = R;
  // function: set pure=false ONLY WIRE
  // function: setby pure=false ONLY WIRE
  // function: get pure=true ONLY WIRE
  sumwrap_uint16_to3 #(.INSTANCE_NAME("regby_inner")) regby_inner(.CLK(CLK), .CE(CE), .process_input({setby_inp,R}), .process_output(regby_inner_process_output));
endmodule

module ChangeRate_uint8_4_1__from8_to2_H1(input CLK, output ready, input reset, input CE, input process_valid, input [255:0] process_input, output [64:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  wire [15:0] phase_GET_OUTPUT;
  wire unnamedbinop12263_readingUSEDMULTIPLEbinop = {(phase_GET_OUTPUT==(16'd0))};
  assign ready = unnamedbinop12263_readingUSEDMULTIPLEbinop;
  reg [63:0] SR_2;
  wire [63:0] unnamedselect12279USEDMULTIPLEselect = ((unnamedbinop12263_readingUSEDMULTIPLEbinop)?(({process_input[63:0]})):(SR_2));
  reg [63:0] unnamedselect12279_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect12279_delay1_validunnamednull0_CECE <= unnamedselect12279USEDMULTIPLEselect; end end
  reg [63:0] SR_1;  always @ (posedge CLK) begin if (process_valid && CE) begin SR_1 <= unnamedselect12279USEDMULTIPLEselect; end end
  reg [63:0] SR_3;
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_2 <= ((unnamedbinop12263_readingUSEDMULTIPLEbinop)?(({process_input[127:64]})):(SR_3)); end end
  reg [63:0] SR_4;
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_3 <= ((unnamedbinop12263_readingUSEDMULTIPLEbinop)?(({process_input[191:128]})):(SR_4)); end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_4 <= ((unnamedbinop12263_readingUSEDMULTIPLEbinop)?(({process_input[255:192]})):(SR_1)); end end
  wire [15:0] phase_SETBY_OUTPUT;
  assign process_output = {(1'd1),unnamedselect12279_delay1_validunnamednull0_CECE};
  // function: ready pure=true delay=0
  // function: reset pure=false delay=0
  // function: process pure=false delay=1
  RegBy_sumwrap_uint16_to3_CEtrue_initnil #(.INSTANCE_NAME("phase")) phase(.CLK(CLK), .set_valid(reset), .CE(CE), .set_inp((16'd0)), .setby_valid(process_valid), .setby_inp((16'd1)), .SETBY_OUTPUT(phase_SETBY_OUTPUT), .GET_OUTPUT(phase_GET_OUTPUT));
endmodule

module WaitOnInput_ChangeRate_uint8_4_1__from8_to2_H1(input CLK, output ready, input reset, input CE, input process_valid, input [256:0] process_input, output [64:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  wire WaitOnInput_inner_ready;
  assign ready = WaitOnInput_inner_ready;
  wire unnamedbinop12385USEDMULTIPLEbinop = {({({(~WaitOnInput_inner_ready)}||(process_input[256]))}&&process_valid)};
  wire [64:0] WaitOnInput_inner_process_output;
  reg unnamedbinop12385_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedbinop12385_delay1_validunnamednull0_CECE <= unnamedbinop12385USEDMULTIPLEbinop; end end
  assign process_output = {{((WaitOnInput_inner_process_output[64])&&unnamedbinop12385_delay1_validunnamednull0_CECE)},(WaitOnInput_inner_process_output[63:0])};
  // function: ready pure=true delay=0
  // function: reset pure=false delay=0
  // function: process pure=false delay=1
  ChangeRate_uint8_4_1__from8_to2_H1 #(.INSTANCE_NAME("WaitOnInput_inner")) WaitOnInput_inner(.CLK(CLK), .ready(WaitOnInput_inner_ready), .reset(reset), .CE(CE), .process_valid(unnamedbinop12385USEDMULTIPLEbinop), .process_input((process_input[255:0])), .process_output(WaitOnInput_inner_process_output));
endmodule

module LiftHandshake_WaitOnInput_ChangeRate_uint8_4_1__from8_to2_H1(input CLK, input ready_downstream, output ready, input reset, input [256:0] process_input, output [64:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire inner_WaitOnInput_ChangeRate_uint8_4_1__from8_to2_H1_ready;
  assign ready = {(inner_WaitOnInput_ChangeRate_uint8_4_1__from8_to2_H1_ready&&ready_downstream)};
  wire unnamedbinop12420USEDMULTIPLEbinop = {(reset||ready_downstream)};
  wire unnamedunary12421USEDMULTIPLEunary = {(~reset)};
  wire [64:0] inner_WaitOnInput_ChangeRate_uint8_4_1__from8_to2_H1_process_output;
  wire validBitDelay_WaitOnInput_ChangeRate_uint8_4_1__from8_to2_H1_pushPop_out;
  wire [64:0] unnamedtuple12431USEDMULTIPLEtuple = {{((inner_WaitOnInput_ChangeRate_uint8_4_1__from8_to2_H1_process_output[64])&&validBitDelay_WaitOnInput_ChangeRate_uint8_4_1__from8_to2_H1_pushPop_out)},(inner_WaitOnInput_ChangeRate_uint8_4_1__from8_to2_H1_process_output[63:0])};
  always @(posedge CLK) begin if({(~{((unnamedtuple12431USEDMULTIPLEtuple[64])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: output valid bit should not be X!",INSTANCE_NAME); end end
  always @(posedge CLK) begin if({(~{((process_input[256])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = unnamedtuple12431USEDMULTIPLEtuple;
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  WaitOnInput_ChangeRate_uint8_4_1__from8_to2_H1 #(.INSTANCE_NAME("inner_WaitOnInput_ChangeRate_uint8_4_1__from8_to2_H1")) inner_WaitOnInput_ChangeRate_uint8_4_1__from8_to2_H1(.CLK(CLK), .ready(inner_WaitOnInput_ChangeRate_uint8_4_1__from8_to2_H1_ready), .reset(reset), .CE(unnamedbinop12420USEDMULTIPLEbinop), .process_valid(unnamedunary12421USEDMULTIPLEunary), .process_input(process_input), .process_output(inner_WaitOnInput_ChangeRate_uint8_4_1__from8_to2_H1_process_output));
  ShiftRegister_1_CEtrue_TY1 #(.INSTANCE_NAME("validBitDelay_WaitOnInput_ChangeRate_uint8_4_1__from8_to2_H1")) validBitDelay_WaitOnInput_ChangeRate_uint8_4_1__from8_to2_H1(.CLK(CLK), .pushPop_valid(unnamedunary12421USEDMULTIPLEunary), .CE(unnamedbinop12420USEDMULTIPLEbinop), .sr_input((1'd1)), .pushPop_out(validBitDelay_WaitOnInput_ChangeRate_uint8_4_1__from8_to2_H1_pushPop_out), .reset(reset));
endmodule

module hsfnfin(input CLK, input ready_downstream, output ready, input reset, input [64:0] process_input, output [64:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire incrate_ready;
  wire O1_ready;
  assign ready = O1_ready;
  wire [256:0] O1_process_output;
  wire [64:0] incrate_process_output;
  assign process_output = incrate_process_output;
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  hsfn #(.INSTANCE_NAME("O1")) O1(.CLK(CLK), .ready_downstream(incrate_ready), .ready(O1_ready), .reset(reset), .process_input(process_input), .process_output(O1_process_output));
  LiftHandshake_WaitOnInput_ChangeRate_uint8_4_1__from8_to2_H1 #(.INSTANCE_NAME("incrate")) incrate(.CLK(CLK), .ready_downstream(ready_downstream), .ready(incrate_ready), .reset(reset), .process_input(O1_process_output), .process_output(incrate_process_output));
endmodule

module Overflow_153600(input CLK, input process_valid, input CE, input [63:0] process_input, output [64:0] process_output, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  reg [63:0] process_input_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_input_delay1_validunnamednull0_CECE <= process_input; end end
  wire [31:0] cnt_GET_OUTPUT;
  reg unnamedbinop12637_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedbinop12637_delay1_validunnamednull0_CECE <= {((cnt_GET_OUTPUT)<((32'd153600)))}; end end
  wire [31:0] cnt_SETBY_OUTPUT;
  assign process_output = {unnamedbinop12637_delay1_validunnamednull0_CECE,process_input_delay1_validunnamednull0_CECE};
  // function: process pure=false delay=1
  // function: reset pure=false delay=0
  RegBy_incif_1uint32_CEtrue_initnil #(.INSTANCE_NAME("cnt")) cnt(.CLK(CLK), .set_valid(reset), .CE(CE), .set_inp((32'd0)), .setby_valid(process_valid), .setby_inp((1'd1)), .SETBY_OUTPUT(cnt_SETBY_OUTPUT), .GET_OUTPUT(cnt_GET_OUTPUT));
endmodule

module LiftDecimate_Overflow_153600(input CLK, output ready, input reset, input CE, input process_valid, input [64:0] process_input, output [64:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  assign ready = (1'd1);
  wire unnamedcast12665USEDMULTIPLEcast = (process_input[64]);
  wire [64:0] LiftDecimate_inner_Overflow_153600_process_output;
  reg [63:0] unnamedcast12668_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast12668_delay1_validunnamednull0_CECE <= (LiftDecimate_inner_Overflow_153600_process_output[63:0]); end end
  reg unnamedcast12665_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast12665_delay1_validunnamednull0_CECE <= unnamedcast12665USEDMULTIPLEcast; end end
  reg unnamedbinop12673_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedbinop12673_delay1_validunnamednull0_CECE <= {((LiftDecimate_inner_Overflow_153600_process_output[64])&&unnamedcast12665_delay1_validunnamednull0_CECE)}; end end
  assign process_output = {unnamedbinop12673_delay1_validunnamednull0_CECE,unnamedcast12668_delay1_validunnamednull0_CECE};
  // function: ready pure=true delay=0
  // function: reset pure=false delay=0
  // function: process pure=false delay=2
  Overflow_153600 #(.INSTANCE_NAME("LiftDecimate_inner_Overflow_153600")) LiftDecimate_inner_Overflow_153600(.CLK(CLK), .process_valid({(unnamedcast12665USEDMULTIPLEcast&&process_valid)}), .CE(CE), .process_input((process_input[63:0])), .process_output(LiftDecimate_inner_Overflow_153600_process_output), .reset(reset));
endmodule

module ShiftRegister_2_CEtrue_TY1(input CLK, input pushPop_valid, input CE, input sr_input, output pushPop_out, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'pushPop'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  reg SR2;
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR1' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR1' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR1' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate12740USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(sr_input):((1'd0)))};
  reg SR1;  always @ (posedge CLK) begin if ((unnamedcallArbitrate12740USEDMULTIPLEcallArbitrate[1]) && CE) begin SR1 <= (unnamedcallArbitrate12740USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR2' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR2' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR2' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate12746USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR1):((1'd0)))};
    always @ (posedge CLK) begin if ((unnamedcallArbitrate12746USEDMULTIPLEcallArbitrate[1]) && CE) begin SR2 <= (unnamedcallArbitrate12746USEDMULTIPLEcallArbitrate[0]); end end
  assign pushPop_out = SR2;
  // function: pushPop pure=false delay=0
  // function: reset pure=false delay=0
endmodule

module LiftHandshake_LiftDecimate_Overflow_153600(input CLK, input ready_downstream, output ready, input reset, input [64:0] process_input, output [64:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire inner_LiftDecimate_Overflow_153600_ready;
  assign ready = {(inner_LiftDecimate_Overflow_153600_ready&&ready_downstream)};
  wire unnamedbinop12710USEDMULTIPLEbinop = {(reset||ready_downstream)};
  wire unnamedunary12711USEDMULTIPLEunary = {(~reset)};
  wire [64:0] inner_LiftDecimate_Overflow_153600_process_output;
  wire validBitDelay_LiftDecimate_Overflow_153600_pushPop_out;
  wire [64:0] unnamedtuple12760USEDMULTIPLEtuple = {{((inner_LiftDecimate_Overflow_153600_process_output[64])&&validBitDelay_LiftDecimate_Overflow_153600_pushPop_out)},(inner_LiftDecimate_Overflow_153600_process_output[63:0])};
  always @(posedge CLK) begin if({(~{((unnamedtuple12760USEDMULTIPLEtuple[64])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: output valid bit should not be X!",INSTANCE_NAME); end end
  always @(posedge CLK) begin if({(~{((process_input[64])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = unnamedtuple12760USEDMULTIPLEtuple;
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  LiftDecimate_Overflow_153600 #(.INSTANCE_NAME("inner_LiftDecimate_Overflow_153600")) inner_LiftDecimate_Overflow_153600(.CLK(CLK), .ready(inner_LiftDecimate_Overflow_153600_ready), .reset(reset), .CE(unnamedbinop12710USEDMULTIPLEbinop), .process_valid(unnamedunary12711USEDMULTIPLEunary), .process_input(process_input), .process_output(inner_LiftDecimate_Overflow_153600_process_output));
  ShiftRegister_2_CEtrue_TY1 #(.INSTANCE_NAME("validBitDelay_LiftDecimate_Overflow_153600")) validBitDelay_LiftDecimate_Overflow_153600(.CLK(CLK), .pushPop_valid(unnamedunary12711USEDMULTIPLEunary), .CE(unnamedbinop12710USEDMULTIPLEbinop), .sr_input((1'd1)), .pushPop_out(validBitDelay_LiftDecimate_Overflow_153600_pushPop_out), .reset(reset));
endmodule

module Underflow_Auint8_4_1__2_1__count153600_cycles154624_toosoonnil_USfalse(input CLK, input ready_downstream, output ready, input reset, input [64:0] process_input, output [64:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  assign ready = ready_downstream;
  wire unnamedbinop13167USEDMULTIPLEbinop = {(ready_downstream||reset)};
  wire [31:0] cycleCount_GET_OUTPUT;
  wire unnamedbinop13166USEDMULTIPLEbinop = {((cycleCount_GET_OUTPUT)>((32'd154624)))};
  wire [31:0] outputCount_GET_OUTPUT;
  wire unnamedcast13160USEDMULTIPLEcast = (process_input[64]);
  wire unnamedunary13186USEDMULTIPLEunary = {(~reset)};
  wire [31:0] outputCount_SETBY_OUTPUT;
  wire [31:0] cycleCount_SETBY_OUTPUT;
  assign process_output = {{({({(unnamedbinop13166USEDMULTIPLEbinop&&{((outputCount_GET_OUTPUT)<((32'd153600)))})}||{({(~unnamedbinop13166USEDMULTIPLEbinop)}&&unnamedcast13160USEDMULTIPLEcast)})}&&unnamedunary13186USEDMULTIPLEunary)},((unnamedbinop13166USEDMULTIPLEbinop)?((64'd3735928559)):((process_input[63:0])))};
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  RegBy_incif_1uint32_CEtrue_initnil #(.INSTANCE_NAME("outputCount")) outputCount(.CLK(CLK), .set_valid(reset), .CE(unnamedbinop13167USEDMULTIPLEbinop), .set_inp((32'd0)), .setby_valid(unnamedunary13186USEDMULTIPLEunary), .setby_inp({(ready_downstream&&{(unnamedcast13160USEDMULTIPLEcast||unnamedbinop13166USEDMULTIPLEbinop)})}), .SETBY_OUTPUT(outputCount_SETBY_OUTPUT), .GET_OUTPUT(outputCount_GET_OUTPUT));
  RegBy_incif_1uint32_CEtrue_initnil #(.INSTANCE_NAME("cycleCount")) cycleCount(.CLK(CLK), .set_valid(reset), .CE(unnamedbinop13167USEDMULTIPLEbinop), .set_inp((32'd0)), .setby_valid(unnamedunary13186USEDMULTIPLEunary), .setby_inp((1'd1)), .SETBY_OUTPUT(cycleCount_SETBY_OUTPUT), .GET_OUTPUT(cycleCount_GET_OUTPUT));
endmodule

module harnessaxi(input CLK, input ready_downstream, output ready, input reset, input [64:0] process_input, output [64:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire underflow_ready;
  wire overflow_ready;
  wire hsfna_ready;
  wire underflow_US_ready;
  assign ready = underflow_US_ready;
  wire [64:0] underflow_US_process_output;
  wire [64:0] hsfna_process_output;
  wire [64:0] overflow_process_output;
  wire [64:0] underflow_process_output;
  assign process_output = underflow_process_output;
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  Underflow_Auint8_8_1__count38400_cycles154624_toosoonnil_UStrue #(.INSTANCE_NAME("underflow_US")) underflow_US(.CLK(CLK), .ready_downstream(hsfna_ready), .ready(underflow_US_ready), .reset(reset), .process_input(process_input), .process_output(underflow_US_process_output));
  hsfnfin #(.INSTANCE_NAME("hsfna")) hsfna(.CLK(CLK), .ready_downstream(overflow_ready), .ready(hsfna_ready), .reset(reset), .process_input(underflow_US_process_output), .process_output(hsfna_process_output));
  LiftHandshake_LiftDecimate_Overflow_153600 #(.INSTANCE_NAME("overflow")) overflow(.CLK(CLK), .ready_downstream(underflow_ready), .ready(overflow_ready), .reset(reset), .process_input(hsfna_process_output), .process_output(overflow_process_output));
  Underflow_Auint8_4_1__2_1__count153600_cycles154624_toosoonnil_USfalse #(.INSTANCE_NAME("underflow")) underflow(.CLK(CLK), .ready_downstream(ready_downstream), .ready(underflow_ready), .reset(reset), .process_input(overflow_process_output), .process_output(underflow_process_output));
endmodule

`timescale 1ps/1ps

module ict106_axilite_conv1 #
  (
   parameter integer C_AXI_ID_WIDTH              = 12,
   parameter integer C_AXI_ADDR_WIDTH            = 32,
   parameter integer C_AXI_DATA_WIDTH            = 32 // CONSTANT
   )
  (
   // System Signals
   input  wire                          ACLK,
   input  wire                          ARESETN,
   input  wire [C_AXI_ID_WIDTH-1:0]     S_AXI_AWID,
   input  wire [C_AXI_ADDR_WIDTH-1:0]   S_AXI_AWADDR,
   input  wire                          S_AXI_AWVALID,
   output wire                          S_AXI_AWREADY,
   input  wire [C_AXI_DATA_WIDTH-1:0]   S_AXI_WDATA,
   input  wire [C_AXI_DATA_WIDTH/8-1:0] S_AXI_WSTRB,
   input  wire                          S_AXI_WVALID,
   output wire                          S_AXI_WREADY,
   output wire [C_AXI_ID_WIDTH-1:0]     S_AXI_BID,
   output wire [2-1:0]                  S_AXI_BRESP,
   output wire                          S_AXI_BVALID,
   input  wire                          S_AXI_BREADY,
   input  wire [C_AXI_ID_WIDTH-1:0]     S_AXI_ARID,
   input  wire [C_AXI_ADDR_WIDTH-1:0]   S_AXI_ARADDR,
   input  wire                          S_AXI_ARVALID,
   output wire                          S_AXI_ARREADY,
   output wire [C_AXI_ID_WIDTH-1:0]     S_AXI_RID,
   output wire [C_AXI_DATA_WIDTH-1:0]   S_AXI_RDATA,
   output wire [2-1:0]                  S_AXI_RRESP,
   output wire                          S_AXI_RLAST,    // Constant =1
   output wire                          S_AXI_RVALID,
   input  wire                          S_AXI_RREADY,
   output wire [C_AXI_ADDR_WIDTH-1:0]   M_AXI_AWADDR,
   output wire                          M_AXI_AWVALID,
   input  wire                          M_AXI_AWREADY,
   output wire [C_AXI_DATA_WIDTH-1:0]   M_AXI_WDATA,
   output wire [C_AXI_DATA_WIDTH/8-1:0] M_AXI_WSTRB,
   output wire                          M_AXI_WVALID,
   input  wire                          M_AXI_WREADY,
   input  wire [2-1:0]                  M_AXI_BRESP,
   input  wire                          M_AXI_BVALID,
   output wire                          M_AXI_BREADY,
   output wire [C_AXI_ADDR_WIDTH-1:0]   M_AXI_ARADDR,
   output wire                          M_AXI_ARVALID,
   input  wire                          M_AXI_ARREADY,
   input  wire [C_AXI_DATA_WIDTH-1:0]   M_AXI_RDATA,
   input  wire [2-1:0]                  M_AXI_RRESP,
   input  wire                          M_AXI_RVALID,
   output wire                          M_AXI_RREADY
  );
  
  wire [31:0] m_axaddr;

  // Arbiter
  reg read_active;
  reg write_active;
  reg busy;

  wire read_req;
  wire write_req;
  wire read_complete;
  wire write_complete;
  
  reg [1:0] areset_d; // Reset delay register
  always @(posedge ACLK) begin
    areset_d <= {areset_d[0], ~ARESETN};
  end
  
  assign read_req  = S_AXI_ARVALID & ~write_active & ~busy & ~|areset_d;
  assign write_req = (S_AXI_AWVALID & ~read_active & ~busy & ~S_AXI_ARVALID & ~|areset_d) | (write_active & ~busy);

  assign read_complete  = M_AXI_RVALID & S_AXI_RREADY;
  assign write_complete = M_AXI_BVALID & S_AXI_BREADY;

  always @(posedge ACLK) begin : arbiter_read_ff
    if (~ARESETN)
      read_active <= 1'b0;
    else if (read_complete)
      read_active <= 1'b0;
    else if (read_req)
      read_active <= 1'b1;
  end

  always @(posedge ACLK) begin : arbiter_write_ff
    if (~ARESETN)
      write_active <= 1'b0;
    else if (write_complete)
      write_active <= 1'b0;
    else if (write_req)
      write_active <= 1'b1;
  end

  always @(posedge ACLK) begin : arbiter_busy_ff
    if (~ARESETN)
      busy <= 1'b0;
    else if (read_complete | write_complete)
      busy <= 1'b0;
    else if ((S_AXI_AWVALID & M_AXI_AWREADY & ~read_req) | (S_AXI_ARVALID & M_AXI_ARREADY & ~write_req))
      busy <= 1'b1;
  end

  assign M_AXI_ARVALID = read_req;
  assign S_AXI_ARREADY = M_AXI_ARREADY & read_req;

  assign M_AXI_AWVALID = write_req;
  assign S_AXI_AWREADY = M_AXI_AWREADY & write_req;

  assign M_AXI_RREADY  = S_AXI_RREADY & read_active;
  assign S_AXI_RVALID  = M_AXI_RVALID & read_active;

  assign M_AXI_BREADY  = S_AXI_BREADY & write_active;
  assign S_AXI_BVALID  = M_AXI_BVALID & write_active;

  // Address multiplexer
  assign m_axaddr = (read_req) ? S_AXI_ARADDR : S_AXI_AWADDR;

  // Id multiplexer and flip-flop
  reg [C_AXI_ID_WIDTH-1:0] s_axid;

  always @(posedge ACLK) begin : axid
    if      (~ARESETN)    s_axid <= {C_AXI_ID_WIDTH{1'b0}};
    else if (read_req)  s_axid <= S_AXI_ARID;
    else if (write_req) s_axid <= S_AXI_AWID;
  end

  assign S_AXI_BID = s_axid;
  assign S_AXI_RID = s_axid;

  assign M_AXI_AWADDR = m_axaddr;
  assign M_AXI_ARADDR = m_axaddr;


  // Feed-through signals
  assign S_AXI_WREADY   = M_AXI_WREADY & ~|areset_d;
  assign S_AXI_BRESP    = M_AXI_BRESP;
  assign S_AXI_RDATA    = M_AXI_RDATA;
  assign S_AXI_RRESP    = M_AXI_RRESP;
  assign S_AXI_RLAST    = 1'b1;

  assign M_AXI_WVALID   = S_AXI_WVALID & ~|areset_d;
  assign M_AXI_WDATA    = S_AXI_WDATA;
  assign M_AXI_WSTRB    = S_AXI_WSTRB;

endmodule

module Conf(
    input ACLK,
    input ARESETN,
    //AXI Inputs
    input [31:0] S_AXI_ARADDR,
    input [11:0] S_AXI_ARID,
    output S_AXI_ARREADY,
    input S_AXI_ARVALID,
    input [31:0] S_AXI_AWADDR,
    input [11:0] S_AXI_AWID,
    output S_AXI_AWREADY,
    input S_AXI_AWVALID,
    output [11:0] S_AXI_BID,
    input S_AXI_BREADY,
    output [1:0] S_AXI_BRESP,
    output S_AXI_BVALID,
    output [31:0] S_AXI_RDATA,
    output [11:0] S_AXI_RID,
    output S_AXI_RLAST,
    input S_AXI_RREADY,
    output [1:0] S_AXI_RRESP,
    output S_AXI_RVALID,
    input [31:0] S_AXI_WDATA,
    output S_AXI_WREADY,
    input [3:0] S_AXI_WSTRB,
    input S_AXI_WVALID,
    
    output CONFIG_VALID,
    input CONFIG_READY,
    output [31:0] CONFIG_CMD,
    output [31:0] CONFIG_SRC,
    output [31:0] CONFIG_DEST,
    output [31:0] CONFIG_LEN,
    output CONFIG_IRQ
    );

    //Convert Input signals to AXI lite, to avoid ID matching
    wire [31:0] LITE_ARADDR;
    wire LITE_ARREADY;
    wire LITE_ARVALID;
    wire [31:0] LITE_AWADDR;
    wire LITE_AWREADY;
    wire LITE_AWVALID;
    wire LITE_BREADY;
    reg [1:0] LITE_BRESP;
    wire LITE_BVALID;
    reg [31:0] LITE_RDATA;
    wire LITE_RREADY;
    reg [1:0] LITE_RRESP;
    wire LITE_RVALID;
    wire [31:0] LITE_WDATA;
    wire LITE_WREADY;
    wire [3:0] LITE_WSTRB;
    wire LITE_WVALID;
    
    ict106_axilite_conv axilite(
    .ACLK(ACLK),
    .ARESETN(ARESETN),
    .S_AXI_ARADDR(S_AXI_ARADDR), 
    .S_AXI_ARID(S_AXI_ARID),  
    .S_AXI_ARREADY(S_AXI_ARREADY), 
    .S_AXI_ARVALID(S_AXI_ARVALID), 
    .S_AXI_AWADDR(S_AXI_AWADDR), 
    .S_AXI_AWID(S_AXI_AWID), 
    .S_AXI_AWREADY(S_AXI_AWREADY), 
    .S_AXI_AWVALID(S_AXI_AWVALID), 
    .S_AXI_BID(S_AXI_BID), 
    .S_AXI_BREADY(S_AXI_BREADY), 
    .S_AXI_BRESP(S_AXI_BRESP), 
    .S_AXI_BVALID(S_AXI_BVALID), 
    .S_AXI_RDATA(S_AXI_RDATA), 
    .S_AXI_RID(S_AXI_RID), 
    .S_AXI_RLAST(S_AXI_RLAST), 
    .S_AXI_RREADY(S_AXI_RREADY), 
    .S_AXI_RRESP(S_AXI_RRESP), 
    .S_AXI_RVALID(S_AXI_RVALID), 
    .S_AXI_WDATA(S_AXI_WDATA), 
    .S_AXI_WREADY(S_AXI_WREADY), 
    .S_AXI_WSTRB(S_AXI_WSTRB), 
    .S_AXI_WVALID(S_AXI_WVALID),
       
    .M_AXI_ARADDR(LITE_ARADDR),
    .M_AXI_ARREADY(LITE_ARREADY),
    .M_AXI_ARVALID(LITE_ARVALID),
    .M_AXI_AWADDR(LITE_AWADDR),
    .M_AXI_AWREADY(LITE_AWREADY),
    .M_AXI_AWVALID(LITE_AWVALID),
    .M_AXI_BREADY(LITE_BREADY),
    .M_AXI_BRESP(LITE_BRESP),
    .M_AXI_BVALID(LITE_BVALID),
    .M_AXI_RDATA(LITE_RDATA),
    .M_AXI_RREADY(LITE_RREADY),
    .M_AXI_RRESP(LITE_RRESP),
    .M_AXI_RVALID(LITE_RVALID),
    .M_AXI_WDATA(LITE_WDATA),
    .M_AXI_WREADY(LITE_WREADY),
    .M_AXI_WSTRB(LITE_WSTRB),
    .M_AXI_WVALID(LITE_WVALID)
  );

parameter NREG = 4;
parameter W = 32;

reg [W-1:0] data[NREG-1:0];

parameter IDLE = 0, RWAIT = 1;
parameter OK = 2'b00, SLVERR = 2'b10;

reg [31:0] counter;

//READS
reg r_state;
wire [1:0] r_select;
assign r_select  = LITE_ARADDR[3:2];
assign ar_good = {LITE_ARADDR[31:4], 2'b00, LITE_ARADDR[1:0]} == 32'h70000000;
assign LITE_ARREADY = (r_state == IDLE);
assign LITE_RVALID = (r_state == RWAIT);
always @(posedge ACLK) begin
    if(ARESETN == 0) begin
        r_state <= IDLE;
    end else case(r_state)
        IDLE: begin
            if(LITE_ARVALID) begin
                LITE_RRESP <= ar_good ? OK : SLVERR;
                LITE_RDATA <= (r_select == 2'b0) ? counter : data[r_select];
                r_state <= RWAIT;
            end
        end
        RWAIT: begin
            if(LITE_RREADY)
                r_state <= IDLE;
        end
    endcase
end 

//WRITES
reg w_state;
reg [1:0] w_select_r;
reg w_wrotedata;
reg w_wroteresp;

wire [1:0] w_select;
assign w_select  = LITE_AWADDR[3:2];
assign aw_good = {LITE_AWADDR[31:4], 2'b00, LITE_AWADDR[1:0]} == 32'h70000000;

assign LITE_AWREADY = (w_state == IDLE);
assign LITE_WREADY = (w_state == RWAIT) && !w_wrotedata;
assign LITE_BVALID = (w_state == RWAIT) && !w_wroteresp;

always @(posedge ACLK) begin
    if(ARESETN == 0) begin
        w_state <= IDLE;
        w_wrotedata <= 0;
        w_wroteresp <= 0;
    end else case(w_state)
        IDLE: begin
            if(LITE_AWVALID) begin
                LITE_BRESP <= aw_good ? OK : SLVERR;
                w_select_r <= w_select;
                w_state <= RWAIT; 
                w_wrotedata <= 0;
                w_wroteresp <= 0;
            end
        end
        RWAIT: begin
            if (LITE_WREADY)
                data[w_select_r] <= LITE_WDATA;
            if((w_wrotedata || LITE_WVALID) && (w_wroteresp || LITE_BREADY)) begin
                w_wrotedata <= 0;
                w_wroteresp <= 0;
                w_state <= IDLE;
            end else if (LITE_WVALID)
                w_wrotedata <= 1;
            else if (LITE_BREADY)
                w_wroteresp <= 1;
        end
    endcase
end

reg v_state;
assign CONFIG_VALID = (v_state == RWAIT);
always @(posedge ACLK) begin
    if (ARESETN == 0)
        v_state <= IDLE;
    else case(v_state)
        IDLE:
            if (LITE_WVALID && LITE_WREADY && w_select_r == 2'b00)
                v_state <= RWAIT;
        RWAIT:
            if (CONFIG_READY)
                v_state <= IDLE;
    endcase
end

assign CONFIG_CMD = data[0];
assign CONFIG_SRC = data[1];
assign CONFIG_DEST = data[2];
assign CONFIG_LEN = data[3];


//how many cycles does the operation take?
always @(posedge ACLK) begin
    if (ARESETN == 0)
        counter <= 0;
    else if (CONFIG_READY && CONFIG_VALID)
        counter <= 0;
    else if (!CONFIG_READY)
        counter <= counter + 1;
end

reg busy;
reg busy_last;
always @(posedge ACLK) begin
    if (ARESETN == 0) begin
        busy <= 0;
        busy_last <= 0;
    end else begin
        if (CONFIG_READY) begin
            busy <= CONFIG_VALID ? 1 : 0;
        end
        busy_last <= busy;
    end
end

assign CONFIG_IRQ = !busy;

endmodule // Conf

module DRAMReader(
    //AXI port
    input ACLK,
    input ARESETN,
    output reg [31:0] M_AXI_ARADDR,
    input M_AXI_ARREADY,
    output  M_AXI_ARVALID,
    input [63:0] M_AXI_RDATA,
    output M_AXI_RREADY,
    input [1:0] M_AXI_RRESP,
    input M_AXI_RVALID,
    input M_AXI_RLAST,
    output [3:0] M_AXI_ARLEN,
    output [1:0] M_AXI_ARSIZE,
    output [1:0] M_AXI_ARBURST,
    
    //Control config
    input CONFIG_VALID,
    output CONFIG_READY,
    input [31:0] CONFIG_START_ADDR,
    input [31:0] CONFIG_NBYTES,
    
    //RAM port
    input DATA_READY_DOWNSTREAM,
    output DATA_VALID,
    output [63:0] DATA
);

assign M_AXI_ARLEN = 4'b1111;
assign M_AXI_ARSIZE = 2'b11;
assign M_AXI_ARBURST = 2'b01;
parameter IDLE = 0, RWAIT = 1;
    
//ADDR logic
reg [31:0] a_count;
reg a_state;  
assign M_AXI_ARVALID = (a_state == RWAIT);
always @(posedge ACLK) begin
    if (ARESETN == 0) begin
        a_state <= IDLE;
        M_AXI_ARADDR <= 0;
        a_count <= 0;
    end else case(a_state)
        IDLE: begin
            if(CONFIG_VALID) begin
                M_AXI_ARADDR <= CONFIG_START_ADDR;
                a_count <= CONFIG_NBYTES[31:7];
                a_state <= RWAIT;
            end
        end
        RWAIT: begin
            if (M_AXI_ARREADY == 1) begin
                if(a_count - 1 == 0)
                    a_state <= IDLE;
                a_count <= a_count - 1;
                M_AXI_ARADDR <= M_AXI_ARADDR + 128; // Bursts are 128 bytes long
            end
        end
    endcase
end
    
//READ logic
reg [31:0] b_count;
reg r_state;
assign M_AXI_RREADY = (r_state == RWAIT) && DATA_READY_DOWNSTREAM;
always @(posedge ACLK) begin
    if (ARESETN == 0) begin
        r_state <= IDLE;
        b_count <= 0;
    end else case(r_state)
        IDLE: begin
            if(CONFIG_VALID) begin
                b_count <= {CONFIG_NBYTES[31:7],7'b0}; // round to nearest 128 bytes
                r_state <= RWAIT;
            end
        end
        RWAIT: begin
            if (M_AXI_RVALID && DATA_READY_DOWNSTREAM) begin
                //use M_AXI_RDATA
                if(b_count - 8 == 0)
                    r_state <= IDLE;
                b_count <= b_count - 8; // each valid cycle the bus provides 8 bytes
            end
        end
    endcase
end

assign DATA = M_AXI_RDATA;
assign DATA_VALID = M_AXI_RVALID && (r_state == RWAIT);
assign CONFIG_READY = (r_state == IDLE) && (a_state == IDLE);

endmodule // DRAMReader

module DRAMWriter(
    //AXI port
    input ACLK,
    input ARESETN,
    output reg [31:0] M_AXI_AWADDR,
    input M_AXI_AWREADY,
    output M_AXI_AWVALID,
    
    output [63:0] M_AXI_WDATA,
    output [7:0] M_AXI_WSTRB,
    input M_AXI_WREADY,
    output M_AXI_WVALID,
    output M_AXI_WLAST,
    
    input [1:0] M_AXI_BRESP,
    input M_AXI_BVALID,
    output M_AXI_BREADY,
    
    output [3:0] M_AXI_AWLEN,
    output [1:0] M_AXI_AWSIZE,
    output [1:0] M_AXI_AWBURST,
    
    //Control config
    input CONFIG_VALID,
    output CONFIG_READY,
    input [31:0] CONFIG_START_ADDR,
    input [31:0] CONFIG_NBYTES,
    
    //RAM port
    input [63:0] DATA,
    output DATA_READY,
    input DATA_VALID

);

assign M_AXI_AWLEN = 4'b1111;
assign M_AXI_AWSIZE = 2'b11;
assign M_AXI_AWBURST = 2'b01;
assign M_AXI_WSTRB = 8'b11111111;

parameter IDLE = 0, RWAIT = 1;
    
//ADDR logic
reg [31:0] a_count;
reg a_state;  
assign M_AXI_AWVALID = (a_state == RWAIT);
always @(posedge ACLK) begin
    if (ARESETN == 0) begin
        a_state <= IDLE;
        M_AXI_AWADDR <= 0;
        a_count <= 0;
    end else case(a_state)
        IDLE: begin
            if(CONFIG_VALID) begin
                M_AXI_AWADDR <= CONFIG_START_ADDR;
                a_count <= CONFIG_NBYTES[31:7];
                a_state <= RWAIT;
            end
        end
        RWAIT: begin
            if (M_AXI_AWREADY == 1) begin
                if(a_count - 1 == 0)
                    a_state <= IDLE;
                a_count <= a_count - 1;
                M_AXI_AWADDR <= M_AXI_AWADDR + 128; 
            end
        end
    endcase
end

//WRITE logic
reg [31:0] b_count;
reg w_state;
always @(posedge ACLK) begin
    if (ARESETN == 0) begin
        w_state <= IDLE;
        b_count <= 0;
    end else case(w_state)
        IDLE: begin
            if(CONFIG_VALID) begin
                b_count <= {CONFIG_NBYTES[31:7],7'b0};
                w_state <= RWAIT;
                last_count <= 4'b1111;
            end
        end
        RWAIT: begin
            if (M_AXI_WREADY && M_AXI_WVALID) begin
                //use M_AXI_WDATA
                if(b_count - 8 == 0) begin
                    w_state <= IDLE;
                end
                last_count <= last_count - 4'b1;
                b_count <= b_count - 8;
            end
        end
    endcase
end

reg [3:0] last_count;
assign M_AXI_WLAST = last_count == 4'b0000;

assign M_AXI_WVALID = (w_state == RWAIT) && DATA_VALID;

assign DATA_READY = (w_state == RWAIT) && M_AXI_WREADY;
   
assign CONFIG_READY = (w_state == IDLE) && (a_state == IDLE);

assign M_AXI_BREADY = 1;

assign M_AXI_WDATA = DATA;

endmodule // DRAMWriter

//-----------------------------------------------------------------------------
// system.v
//-----------------------------------------------------------------------------

// The axi bus expects the number of valid data items to exactly match the # of addresses we send.
// This module checks for underflow (too few valid data items). If there are too few, it inserts DEADBEEFs to make it correct.
// lengthOutput is in bytes
module UnderflowShim(input CLK, input RST, input [31:0] lengthOutput, input [63:0] inp, input inp_valid, output [63:0] out, output out_valid);
   parameter WAIT_CYCLES = 2048;
   
   reg [31:0] outCnt;
   reg [31:0] outLen;

   reg        fixupMode;
   reg [31:0]  outClks = 0;
   
   
   always@(posedge CLK) begin
     if (RST) begin 
        outCnt <= 32'd0;
        outLen <= lengthOutput;
        fixupMode <= 1'b0;
        outClks <= 32'd0;
     end else begin
        outClks <= outClks + 32'd1;
        
        if(inp_valid || fixupMode) begin outCnt <= outCnt+32'd8; end // AXI does 8 bytes per clock
        if(outClks > WAIT_CYCLES) begin fixupMode <= 1'b1; end
     end
   end

   assign out = (fixupMode)?(64'hDEAD):(inp);
   assign out_valid = (RST)?(1'b0):((fixupMode)?(outCnt<outLen):(inp_valid));
endmodule

module stage
  (
    inout [53:0] MIO,
    inout PS_SRSTB,
    inout PS_CLK,
    inout PS_PORB,
    inout DDR_Clk,
    inout DDR_Clk_n,
    inout DDR_CKE,
    inout DDR_CS_n,
    inout DDR_RAS_n,
    inout DDR_CAS_n,
    output DDR_WEB,
    inout [2:0] DDR_BankAddr,
    inout [14:0] DDR_Addr,
    inout DDR_ODT,
    inout DDR_DRSTB,
    inout [31:0] DDR_DQ,
    inout [3:0] DDR_DM,
    inout [3:0] DDR_DQS,
    inout [3:0] DDR_DQS_n,
    inout DDR_VRN,
    inout DDR_VRP,
    output [7:0] LED
  );

  wire [3:0] fclk;
  wire [3:0] fclkresetn;
  wire FCLK0;
  BUFG bufg(.I(fclk[0]),.O(FCLK0));
  assign ARESETN = fclkresetn[0];
  
  
    wire [31:0] PS7_ARADDR;
    wire [11:0] PS7_ARID;
    wire [2:0] PS7_ARPROT;
    wire PS7_ARREADY;
    wire PS7_ARVALID;
    wire [31:0] PS7_AWADDR;
    wire [11:0] PS7_AWID;
    wire [2:0] PS7_AWPROT;
    wire PS7_AWREADY;
    wire PS7_AWVALID;
    wire [11:0] PS7_BID;
    wire PS7_BREADY;
    wire [1:0] PS7_BRESP;
    wire PS7_BVALID;
    wire [31:0] PS7_RDATA;
    wire [11:0] PS7_RID;
    wire PS7_RLAST;
    wire PS7_RREADY;
    wire [1:0] PS7_RRESP;
    wire PS7_RVALID;
    wire [31:0] PS7_WDATA;
    wire PS7_WREADY;
    wire [3:0] PS7_WSTRB;
    wire PS7_WVALID;

    wire [31:0] M_AXI_ARADDR;
    wire M_AXI_ARREADY;
    wire  M_AXI_ARVALID;
    wire [31:0] M_AXI_AWADDR;
    wire M_AXI_AWREADY;
    wire  M_AXI_AWVALID;
    wire  M_AXI_BREADY;
    wire [1:0] M_AXI_BRESP;
    wire M_AXI_BVALID;
    wire [63:0] M_AXI_RDATA;
    wire M_AXI_RREADY;
    wire [1:0] M_AXI_RRESP;
    wire M_AXI_RVALID;
    wire [63:0] M_AXI_WDATA;
    wire M_AXI_WREADY;
    wire [7:0] M_AXI_WSTRB;
    wire M_AXI_WVALID;
    wire M_AXI_RLAST;
    wire M_AXI_WLAST;
    
    wire [3:0] M_AXI_ARLEN;
    wire [1:0] M_AXI_ARSIZE;
    wire [1:0] M_AXI_ARBURST;
    
    wire [3:0] M_AXI_AWLEN;
    wire [1:0] M_AXI_AWSIZE;
    wire [1:0] M_AXI_AWBURST;
    
    wire CONFIG_VALID;
    wire [31:0] CONFIG_CMD;
    wire [31:0] CONFIG_SRC;
    wire [31:0] CONFIG_DEST;
    wire [31:0] CONFIG_LEN;
    wire CONFIG_IRQ;
  
    wire READER_READY;
    wire WRITER_READY;
    
    assign CONFIG_READY = READER_READY && WRITER_READY;
    
    Conf conf(
    .ACLK(FCLK0),
    .ARESETN(ARESETN),
    .S_AXI_ARADDR(PS7_ARADDR), 
    .S_AXI_ARID(PS7_ARID),  
    .S_AXI_ARREADY(PS7_ARREADY), 
    .S_AXI_ARVALID(PS7_ARVALID), 
    .S_AXI_AWADDR(PS7_AWADDR), 
    .S_AXI_AWID(PS7_AWID), 
    .S_AXI_AWREADY(PS7_AWREADY), 
    .S_AXI_AWVALID(PS7_AWVALID), 
    .S_AXI_BID(PS7_BID), 
    .S_AXI_BREADY(PS7_BREADY), 
    .S_AXI_BRESP(PS7_BRESP), 
    .S_AXI_BVALID(PS7_BVALID), 
    .S_AXI_RDATA(PS7_RDATA), 
    .S_AXI_RID(PS7_RID), 
    .S_AXI_RLAST(PS7_RLAST), 
    .S_AXI_RREADY(PS7_RREADY), 
    .S_AXI_RRESP(PS7_RRESP), 
    .S_AXI_RVALID(PS7_RVALID), 
    .S_AXI_WDATA(PS7_WDATA), 
    .S_AXI_WREADY(PS7_WREADY), 
    .S_AXI_WSTRB(PS7_WSTRB), 
    .S_AXI_WVALID(PS7_WVALID),
    .CONFIG_VALID(CONFIG_VALID),
    .CONFIG_READY(CONFIG_READY),
    .CONFIG_CMD(CONFIG_CMD),
    .CONFIG_SRC(CONFIG_SRC),
    .CONFIG_DEST(CONFIG_DEST),
    .CONFIG_LEN(CONFIG_LEN),
    .CONFIG_IRQ(CONFIG_IRQ));

   // lengthInput/lengthOutput are in bytes
   wire [31:0] lengthInput;
   assign lengthInput = {4'b0000,CONFIG_LEN[27:0]};
   wire [31:0] lengthOutput;
   assign lengthOutput = (CONFIG_LEN[27:0] << 8'd8) >> CONFIG_LEN[31:28];

   reg [31:0]  clkcnt = 0;
//   assign LED = clkcnt[20:13];
   assign  LED = clkcnt[28:21];
   
  always @(posedge FCLK0) begin
//    if(ARESETN == 0)
//        LED <= 0;
//    else if(CONFIG_VALID)
//        LED <= {CONFIG_CMD[1:0],CONFIG_SRC[2:0],CONFIG_DEST[2:0]};
     clkcnt <= clkcnt+1;

  end

  wire [63:0] pipelineInput;
  wire       pipelineInputValid;
   
  wire [64:0] pipelineOutputPacked;
  wire [63:0] pipelineOutput;
  assign pipelineOutput = pipelineOutputPacked[63:0];   
  wire pipelineOutputValid;
  assign pipelineOutputValid = pipelineOutputPacked[64];
   
  wire       pipelineReady;
  wire      downstreamReady;

  
    
  harnessaxi  #(.INPUT_COUNT(38400),.OUTPUT_COUNT(153600)) pipeline(.CLK(FCLK0),.reset(CONFIG_READY),.ready(pipelineReady),.ready_downstream(downstreamReady),.process_input({pipelineInputValid,pipelineInput}),.process_output(pipelineOutputPacked));

//   UnderflowShim #(.WAIT_CYCLES(39424)) OS(.CLK(FCLK0),.RST(CONFIG_READY),.lengthOutput(lengthOutput),.inp(pipelineOutputPacked[63:0]),.inp_valid(pipelineOutputPacked[64]),.out(pipelineOutput),.out_valid(pipelineOutputValid));
   
  DRAMReader reader(
    .ACLK(FCLK0),
    .ARESETN(ARESETN),
    .M_AXI_ARADDR(M_AXI_ARADDR),
    .M_AXI_ARREADY(M_AXI_ARREADY),
    .M_AXI_ARVALID(M_AXI_ARVALID),
    .M_AXI_RDATA(M_AXI_RDATA),
    .M_AXI_RREADY(M_AXI_RREADY),
    .M_AXI_RRESP(M_AXI_RRESP),
    .M_AXI_RVALID(M_AXI_RVALID),
    .M_AXI_RLAST(M_AXI_RLAST),
    .M_AXI_ARLEN(M_AXI_ARLEN),
    .M_AXI_ARSIZE(M_AXI_ARSIZE),
    .M_AXI_ARBURST(M_AXI_ARBURST),
    
    .CONFIG_VALID(CONFIG_VALID),
    .CONFIG_READY(READER_READY),
    .CONFIG_START_ADDR(CONFIG_SRC),
    .CONFIG_NBYTES(307200),

    .DATA_READY_DOWNSTREAM(pipelineReady),
    .DATA_VALID(pipelineInputValid),
    .DATA(pipelineInput)
  );
  
  DRAMWriter writer(
    .ACLK(FCLK0),
    .ARESETN(ARESETN),
    .M_AXI_AWADDR(M_AXI_AWADDR),
    .M_AXI_AWREADY(M_AXI_AWREADY),
    .M_AXI_AWVALID(M_AXI_AWVALID),
    .M_AXI_WDATA(M_AXI_WDATA),
    .M_AXI_WREADY(M_AXI_WREADY),
    .M_AXI_WVALID(M_AXI_WVALID),
    .M_AXI_WLAST(M_AXI_WLAST),
    .M_AXI_WSTRB(M_AXI_WSTRB),
    
    .M_AXI_BRESP(M_AXI_BRESP),
    .M_AXI_BREADY(M_AXI_BREADY),
    .M_AXI_BVALID(M_AXI_BVALID),
    
    .M_AXI_AWLEN(M_AXI_AWLEN),
    .M_AXI_AWSIZE(M_AXI_AWSIZE),
    .M_AXI_AWBURST(M_AXI_AWBURST),
    
    .CONFIG_VALID(CONFIG_VALID),
    .CONFIG_READY(WRITER_READY),
    .CONFIG_START_ADDR(CONFIG_DEST),
    .CONFIG_NBYTES(1228800),

    .DATA_READY(downstreamReady),
    .DATA_VALID(pipelineOutputValid),
    .DATA(pipelineOutput)
  );

  PS7 ps7_0(
    .DMA0DATYPE(), 	// out std_logic_vector(1 downto 0);
    .DMA0DAVALID(), 	// out std_ulogic;
    .DMA0DRREADY(), 	// out std_ulogic;
    .DMA0RSTN(), 	// out std_ulogic;
    .DMA1DATYPE(), 	// out std_logic_vector(1 downto 0);
    .DMA1DAVALID(), 	// out std_ulogic;
    .DMA1DRREADY(), 	// out std_ulogic;
    .DMA1RSTN(), 	// out std_ulogic;
    .DMA2DATYPE(), 	// out std_logic_vector(1 downto 0);
    .DMA2DAVALID(), 	// out std_ulogic;
    .DMA2DRREADY(), 	// out std_ulogic;
    .DMA2RSTN(), 	// out std_ulogic;
    .DMA3DATYPE(), 	// out std_logic_vector(1 downto 0);
    .DMA3DAVALID(), 	// out std_ulogic;
    .DMA3DRREADY(), 	// out std_ulogic;
    .DMA3RSTN(), 	// out std_ulogic;
    .EMIOCAN0PHYTX(), 	// out std_ulogic;
    .EMIOCAN1PHYTX(), 	// out std_ulogic;
    .EMIOENET0GMIITXD(), 	// out std_logic_vector(7 downto 0);
    .EMIOENET0GMIITXEN(), 	// out std_ulogic;
    .EMIOENET0GMIITXER(), 	// out std_ulogic;
    .EMIOENET0MDIOMDC(), 	// out std_ulogic;
    .EMIOENET0MDIOO(), 	// out std_ulogic;
    .EMIOENET0MDIOTN(), 	// out std_ulogic;
    .EMIOENET0PTPDELAYREQRX(), 	// out std_ulogic;
    .EMIOENET0PTPDELAYREQTX(), 	// out std_ulogic;
    .EMIOENET0PTPPDELAYREQRX(), 	// out std_ulogic;
    .EMIOENET0PTPPDELAYREQTX(), 	// out std_ulogic;
    .EMIOENET0PTPPDELAYRESPRX(), 	// out std_ulogic;
    .EMIOENET0PTPPDELAYRESPTX(), 	// out std_ulogic;
    .EMIOENET0PTPSYNCFRAMERX(), 	// out std_ulogic;
    .EMIOENET0PTPSYNCFRAMETX(), 	// out std_ulogic;
    .EMIOENET0SOFRX(), 	// out std_ulogic;
    .EMIOENET0SOFTX(), 	// out std_ulogic;
    .EMIOENET1GMIITXD(), 	// out std_logic_vector(7 downto 0);
    .EMIOENET1GMIITXEN(), 	// out std_ulogic;
    .EMIOENET1GMIITXER(), 	// out std_ulogic;
    .EMIOENET1MDIOMDC(), 	// out std_ulogic;
    .EMIOENET1MDIOO(), 	// out std_ulogic;
    .EMIOENET1MDIOTN(), 	// out std_ulogic;
    .EMIOENET1PTPDELAYREQRX(), 	// out std_ulogic;
    .EMIOENET1PTPDELAYREQTX(), 	// out std_ulogic;
    .EMIOENET1PTPPDELAYREQRX(), 	// out std_ulogic;
    .EMIOENET1PTPPDELAYREQTX(), 	// out std_ulogic;
    .EMIOENET1PTPPDELAYRESPRX(), 	// out std_ulogic;
    .EMIOENET1PTPPDELAYRESPTX(), 	// out std_ulogic;
    .EMIOENET1PTPSYNCFRAMERX(), 	// out std_ulogic;
    .EMIOENET1PTPSYNCFRAMETX(), 	// out std_ulogic;
    .EMIOENET1SOFRX(), 	// out std_ulogic;
    .EMIOENET1SOFTX(), 	// out std_ulogic;
    .EMIOGPIOO(), 	 // out std_logic_vector(63 downto 0);
    .EMIOGPIOTN(),  // out std_logic_vector(63 downto 0);
    .EMIOI2C0SCLO(), 	 // out std_ulogic;
    .EMIOI2C0SCLTN(),  // out std_ulogic;
    .EMIOI2C0SDAO(), 	 // out std_ulogic;
    .EMIOI2C0SDATN(),  // out std_ulogic;
    .EMIOI2C1SCLO(), 	 // out std_ulogic;
    .EMIOI2C1SCLTN(),  // out std_ulogic;
    .EMIOI2C1SDAO(), 	 // out std_ulogic;
    .EMIOI2C1SDATN(),  // out std_ulogic;
    .EMIOPJTAGTDO(), 	// out std_ulogic;
    .EMIOPJTAGTDTN(), 	// out std_ulogic;
    .EMIOSDIO0BUSPOW(), 	// out std_ulogic;
    .EMIOSDIO0BUSVOLT(), 	// out std_logic_vector(2 downto 0);
    .EMIOSDIO0CLK(), 	// out std_ulogic;
    .EMIOSDIO0CMDO(), 	// out std_ulogic;
    .EMIOSDIO0CMDTN(), 	// out std_ulogic;
    .EMIOSDIO0DATAO(), 	// out std_logic_vector(3 downto 0);
    .EMIOSDIO0DATATN(), 	// out std_logic_vector(3 downto 0);
    .EMIOSDIO0LED(), 	// out std_ulogic;
    .EMIOSDIO1BUSPOW(), 	// out std_ulogic;
    .EMIOSDIO1BUSVOLT(), 	// out std_logic_vector(2 downto 0);
    .EMIOSDIO1CLK(), 	// out std_ulogic;
    .EMIOSDIO1CMDO(), 	// out std_ulogic;
    .EMIOSDIO1CMDTN(), 	// out std_ulogic;
    .EMIOSDIO1DATAO(), 	// out std_logic_vector(3 downto 0);
    .EMIOSDIO1DATATN(), 	// out std_logic_vector(3 downto 0);
    .EMIOSDIO1LED(), 	// out std_ulogic;
    .EMIOSPI0MO(), 	// out std_ulogic;
    .EMIOSPI0MOTN(), 	// out std_ulogic;
    .EMIOSPI0SCLKO(), 	// out std_ulogic;
    .EMIOSPI0SCLKTN(), 	// out std_ulogic;
    .EMIOSPI0SO(), 	// out std_ulogic;
    .EMIOSPI0SSNTN(), 	// out std_ulogic;
    .EMIOSPI0SSON(), 	// out std_logic_vector(2 downto 0);
    .EMIOSPI0STN(), 	// out std_ulogic;
    .EMIOSPI1MO(), 	// out std_ulogic;
    .EMIOSPI1MOTN(), 	// out std_ulogic;
    .EMIOSPI1SCLKO(), 	// out std_ulogic;
    .EMIOSPI1SCLKTN(), 	// out std_ulogic;
    .EMIOSPI1SO(), 	// out std_ulogic;
    .EMIOSPI1SSNTN(), 	// out std_ulogic;
    .EMIOSPI1SSON(), 	// out std_logic_vector(2 downto 0);
    .EMIOSPI1STN(), 	// out std_ulogic;
    .EMIOTRACECTL(), 	// out std_ulogic;
    .EMIOTRACEDATA(), 	// out std_logic_vector(31 downto 0);
    .EMIOTTC0WAVEO(), 	// out std_logic_vector(2 downto 0);
    .EMIOTTC1WAVEO(), 	// out std_logic_vector(2 downto 0);
    .EMIOUART0DTRN(), 	// out std_ulogic;
    .EMIOUART0RTSN(), 	// out std_ulogic;
    .EMIOUART0TX(), 	// out std_ulogic;
    .EMIOUART1DTRN(), 	// out std_ulogic;
    .EMIOUART1RTSN(), 	// out std_ulogic;
    .EMIOUART1TX(), 	// out std_ulogic;
    .EMIOUSB0PORTINDCTL(), 	// out std_logic_vector(1 downto 0);
    .EMIOUSB0VBUSPWRSELECT(), 	// out std_ulogic;
    .EMIOUSB1PORTINDCTL(), 	// out std_logic_vector(1 downto 0);
    .EMIOUSB1VBUSPWRSELECT(), 	// out std_ulogic;
    .EMIOWDTRSTO(), 	// out std_ulogic;
    .EVENTEVENTO(), 	// out std_ulogic;
    .EVENTSTANDBYWFE(), 	// out std_logic_vector(1 downto 0);
    .EVENTSTANDBYWFI(), 	// out std_logic_vector(1 downto 0);
    .FCLKCLK(fclk), 	 // out std_logic_vector(3 downto 0);
    .FCLKRESETN(fclkresetn), 	// out std_logic_vector(3 downto 0);
    .FTMTF2PTRIGACK(), 	// out std_logic_vector(3 downto 0);
    .FTMTP2FDEBUG(), 	// out std_logic_vector(31 downto 0);
    .FTMTP2FTRIG(), 	// out std_logic_vector(3 downto 0);
    .IRQP2F(), 	// out std_logic_vector(28 downto 0);
    
    .MAXIGP0ACLK(FCLK0), 	// in std_ulogic;
    .MAXIGP0ARADDR(PS7_ARADDR),  // out std_logic_vector(31 downto 0);
    .MAXIGP0ARBURST(),  // out std_logic_vector(1 downto 0);
    .MAXIGP0ARCACHE(),  // out std_logic_vector(3 downto 0);
    .MAXIGP0ARESETN(),  // out std_ulogic;
    .MAXIGP0ARID(PS7_ARID), 	 // out std_logic_vector(11 downto 0);
    .MAXIGP0ARLEN(),  // out std_logic_vector(3 downto 0);
    .MAXIGP0ARLOCK(),  // out std_logic_vector(1 downto 0);
    .MAXIGP0ARPROT(),  // out std_logic_vector(2 downto 0);
    .MAXIGP0ARQOS(),  // out std_logic_vector(3 downto 0);
    .MAXIGP0ARREADY(PS7_ARREADY), // in std_ulogic;
    .MAXIGP0ARSIZE(),  // out std_logic_vector(1 downto 0);
    .MAXIGP0ARVALID(PS7_ARVALID),  // out std_ulogic;
    .MAXIGP0AWADDR(PS7_AWADDR),  // out std_logic_vector(31 downto 0);
    .MAXIGP0AWBURST(),  // out std_logic_vector(1 downto 0);
    .MAXIGP0AWCACHE(),  // out std_logic_vector(3 downto 0);
    .MAXIGP0AWID(PS7_AWID), 	 // out std_logic_vector(11 downto 0);
    .MAXIGP0AWLEN(),  // out std_logic_vector(3 downto 0);
    .MAXIGP0AWLOCK(),  // out std_logic_vector(1 downto 0);
    .MAXIGP0AWPROT(),  // out std_logic_vector(2 downto 0);
    .MAXIGP0AWQOS(),  // out std_logic_vector(3 downto 0);
    .MAXIGP0AWREADY(PS7_AWREADY), // in std_ulogic;
    .MAXIGP0AWSIZE(),  // out std_logic_vector(1 downto 0);
    .MAXIGP0AWVALID(PS7_AWVALID),  // out std_ulogic;
    .MAXIGP0BID(PS7_BID), 	// in std_logic_vector(11 downto 0);
    .MAXIGP0BREADY(PS7_BREADY),  // out std_ulogic;
    .MAXIGP0BRESP(PS7_BRESP), // in std_logic_vector(1 downto 0);
    .MAXIGP0BVALID(PS7_BVALID), // in std_ulogic;
    .MAXIGP0RDATA(PS7_RDATA), // in std_logic_vector(31 downto 0);
    .MAXIGP0RID(PS7_RID), 	// in std_logic_vector(11 downto 0);
    .MAXIGP0RLAST(PS7_RLAST), // in std_ulogic;
    .MAXIGP0RREADY(PS7_RREADY),  // out std_ulogic;
    .MAXIGP0RRESP(PS7_RRESP), // in std_logic_vector(1 downto 0);    
    .MAXIGP0RVALID(PS7_RVALID), // in std_ulogic;
    .MAXIGP0WDATA(PS7_WDATA),  // out std_logic_vector(31 downto 0);
    .MAXIGP0WID(), 	 // out std_logic_vector(11 downto 0);
    .MAXIGP0WLAST(),  // out std_ulogic;
    .MAXIGP0WREADY(PS7_WREADY), // in std_ulogic;
    .MAXIGP0WSTRB(PS7_WSTRB),  // out std_logic_vector(3 downto 0);
    .MAXIGP0WVALID(PS7_WVALID),  // out std_ulogic;
    
    .MAXIGP1ARADDR(),  // out std_logic_vector(31 downto 0);
    .MAXIGP1ARBURST(),  // out std_logic_vector(1 downto 0);
    .MAXIGP1ARCACHE(),  // out std_logic_vector(3 downto 0);
    .MAXIGP1ARESETN(),  // out std_ulogic;
    .MAXIGP1ARID(), 	 // out std_logic_vector(11 downto 0);
    .MAXIGP1ARLEN(),  // out std_logic_vector(3 downto 0);
    .MAXIGP1ARLOCK(),  // out std_logic_vector(1 downto 0);
    .MAXIGP1ARPROT(),  // out std_logic_vector(2 downto 0);
    .MAXIGP1ARQOS(),  // out std_logic_vector(3 downto 0);
    .MAXIGP1ARSIZE(),  // out std_logic_vector(1 downto 0);
    .MAXIGP1ARVALID(),  // out std_ulogic;
    .MAXIGP1AWADDR(),  // out std_logic_vector(31 downto 0);
    .MAXIGP1AWBURST(),  // out std_logic_vector(1 downto 0);
    .MAXIGP1AWCACHE(),  // out std_logic_vector(3 downto 0);
    .MAXIGP1AWID(), 	 // out std_logic_vector(11 downto 0);
    .MAXIGP1AWLEN(),  // out std_logic_vector(3 downto 0);
    .MAXIGP1AWLOCK(),  // out std_logic_vector(1 downto 0);
    .MAXIGP1AWPROT(),  // out std_logic_vector(2 downto 0);
    .MAXIGP1AWQOS(),  // out std_logic_vector(3 downto 0);
    .MAXIGP1AWSIZE(),  // out std_logic_vector(1 downto 0);
    .MAXIGP1AWVALID(),  // out std_ulogic;
    .MAXIGP1BREADY(),  // out std_ulogic;
    .MAXIGP1RREADY(),  // out std_ulogic;
    .MAXIGP1WDATA(),  // out std_logic_vector(31 downto 0);
    .MAXIGP1WID(), 	 // out std_logic_vector(11 downto 0);
    .MAXIGP1WLAST(),  // out std_ulogic;
    .MAXIGP1WSTRB(),  // out std_logic_vector(3 downto 0);
    .MAXIGP1WVALID(),  // out std_ulogic;
    .SAXIGP0ARESETN(), 	// out std_ulogic;
    .SAXIGP0ARREADY(), 	// out std_ulogic;
    .SAXIGP0AWREADY(), 	// out std_ulogic;
    .SAXIGP0BID(), 	// out std_logic_vector(5 downto 0);
    .SAXIGP0BRESP(), 	// out std_logic_vector(1 downto 0);
    .SAXIGP0BVALID(), 	// out std_ulogic;
    .SAXIGP0RDATA(), 	// out std_logic_vector(31 downto 0);
    .SAXIGP0RID(), 	// out std_logic_vector(5 downto 0);
    .SAXIGP0RLAST(), 	// out std_ulogic;
    .SAXIGP0RRESP(), 	// out std_logic_vector(1 downto 0);
    .SAXIGP0RVALID(), 	// out std_ulogic;
    .SAXIGP0WREADY(), 	// out std_ulogic;
    .SAXIGP1ARESETN(), 	// out std_ulogic;
    .SAXIGP1ARREADY(), 	// out std_ulogic;
    .SAXIGP1AWREADY(), 	// out std_ulogic;
    .SAXIGP1BID(), 	// out std_logic_vector(5 downto 0);
    .SAXIGP1BRESP(), 	// out std_logic_vector(1 downto 0);
    .SAXIGP1BVALID(), 	// out std_ulogic;
    .SAXIGP1RDATA(), 	// out std_logic_vector(31 downto 0);
    .SAXIGP1RID(), 	// out std_logic_vector(5 downto 0);
    .SAXIGP1RLAST(), 	// out std_ulogic;
    .SAXIGP1RRESP(), 	// out std_logic_vector(1 downto 0);
    .SAXIGP1RVALID(), 	// out std_ulogic;
    .SAXIGP1WREADY(), 	// out std_ulogic;
    
    
    
    .SAXIHP0ACLK(1'b0), 		// in std_ulogic;
    .SAXIHP0ARADDR(32'b0),	// in std_logic_vector(31 downto 0);
    .SAXIHP0ARBURST(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIHP0ARCACHE(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIHP0ARESETN(), 	// out std_ulogic;
    .SAXIHP0ARID(6'b0),	// in std_logic_vector(2 downto 0);
    .SAXIHP0ARLEN(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIHP0ARLOCK(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIHP0ARPROT(3'b0),	// in std_logic_vector(2 downto 0);
    .SAXIHP0ARQOS(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIHP0ARREADY(), 	// out std_ulogic;
    .SAXIHP0ARSIZE(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIHP0ARVALID(1'b0), 		// in std_ulogic;
    .SAXIHP0AWADDR(32'b0),	// in std_logic_vector(31 downto 0);
    .SAXIHP0AWBURST(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIHP0AWCACHE(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIHP0AWID(6'b0),	// in std_logic_vector(2 downto 0);
    .SAXIHP0AWLEN(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIHP0AWLOCK(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIHP0AWPROT(3'b0),	// in std_logic_vector(2 downto 0);
    .SAXIHP0AWQOS(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIHP0AWREADY(), 	// out std_ulogic;
    .SAXIHP0AWSIZE(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIHP0AWVALID(1'b0), 		// in std_ulogic;
    .SAXIHP0BID(), 	// out std_logic_vector(2 downto 0);
    .SAXIHP0BREADY(1'b0), 		// in std_ulogic;
    .SAXIHP0BRESP(), 	// out std_logic_vector(1 downto 0);
    .SAXIHP0BVALID(), 	// out std_ulogic;
    .SAXIHP0RDATA(), 	// out std_logic_vector(63 downto 0);
    .SAXIHP0RID(), 	// out std_logic_vector(2 downto 0);
    .SAXIHP0RLAST(), 	// out std_ulogic;
    .SAXIHP0RREADY(1'b0), 		// in std_ulogic;
    .SAXIHP0RRESP(), 	// out std_logic_vector(1 downto 0);
    .SAXIHP0RVALID(), 	// out std_ulogic;
    .SAXIHP0WDATA(64'b0),	// in std_logic_vector(63 downto 0);
    .SAXIHP0WID(6'b0),	// in std_logic_vector(2 downto 0);
    .SAXIHP0WLAST(1'b0), 		// in std_ulogic;
    .SAXIHP0WREADY(), 	// out std_ulogic;
    .SAXIHP0WSTRB(8'b0),	// in std_logic_vector(7 downto 0);
    .SAXIHP0WVALID(1'b0), 		// in std_ulogic;
    
    .SAXIACPARUSER(5'b0),	// in std_logic_vector(4 downto 0);
    .SAXIACPAWUSER(5'b0),	// in std_logic_vector(4 downto 0);
    
    .SAXIACPACLK(FCLK0), 	// in std_ulogic;
    .SAXIACPARADDR(M_AXI_ARADDR),
    .SAXIACPARBURST(M_AXI_ARBURST), // in std_logic_vector(1 downto 0);
    .SAXIACPARCACHE(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIACPARESETN(),  // out std_ulogic;
    .SAXIACPARID(3'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIACPARLEN(M_AXI_ARLEN), // in std_logic_vector(3 downto 0);
    .SAXIACPARLOCK(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIACPARPROT(3'b0), // in std_logic_vector(2 downto 0);
    .SAXIACPARQOS(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIACPARREADY(M_AXI_ARREADY),
    .SAXIACPARSIZE(M_AXI_ARSIZE), // in std_logic_vector(1 downto 0);
    .SAXIACPARVALID(M_AXI_ARVALID),
    .SAXIACPAWADDR(M_AXI_AWADDR),
    .SAXIACPAWBURST(M_AXI_AWBURST), // in std_logic_vector(1 downto 0);
    .SAXIACPAWCACHE(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIACPAWID(3'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIACPAWLEN(M_AXI_AWLEN), // in std_logic_vector(3 downto 0);
    .SAXIACPAWLOCK(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIACPAWPROT(3'b0), // in std_logic_vector(2 downto 0);
    .SAXIACPAWQOS(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIACPAWREADY(M_AXI_AWREADY),
    .SAXIACPAWSIZE(M_AXI_AWSIZE), // in std_logic_vector(1 downto 0);
    .SAXIACPAWVALID(M_AXI_AWVALID),
    .SAXIACPBID(), 	 // out std_logic_vector(5 downto 0);
    .SAXIACPBREADY(M_AXI_BREADY),
    .SAXIACPBRESP(M_AXI_BRESP),
    .SAXIACPBVALID(M_AXI_BVALID),
    .SAXIACPRDATA(M_AXI_RDATA),
    .SAXIACPRID(), 	 // out std_logic_vector(5 downto 0);
    .SAXIACPRLAST(M_AXI_RLAST),  // out std_ulogic;
    .SAXIACPRREADY(M_AXI_RREADY),
    .SAXIACPRRESP(M_AXI_RRESP),
    .SAXIACPRVALID(M_AXI_RVALID),
    .SAXIACPWDATA(M_AXI_WDATA),
    .SAXIACPWID(3'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIACPWLAST(M_AXI_WLAST), // in std_ulogic;
    .SAXIACPWREADY(M_AXI_WREADY),
    .SAXIACPWSTRB(M_AXI_WSTRB),
    .SAXIACPWVALID(M_AXI_WVALID),
    
    .SAXIHP0RDISSUECAP1EN(1'b0), 		// in std_ulogic;
    .SAXIHP0WRISSUECAP1EN(1'b0), 		// in std_ulogic;
    .SAXIHP0RACOUNT(),  // out std_logic_vector(2 downto 0);
    .SAXIHP0RCOUNT(),  // out std_logic_vector(7 downto 0);
    .SAXIHP0WACOUNT(),  // out std_logic_vector(5 downto 0);
    .SAXIHP0WCOUNT(),  // out std_logic_vector(7 downto 0);
    
    .SAXIHP1ARESETN(),  // out std_ulogic;
    .SAXIHP1ARREADY(),  // out std_ulogic;
    .SAXIHP1AWREADY(),  // out std_ulogic;
    .SAXIHP1BID(), 	 // out std_logic_vector(5 downto 0);
    .SAXIHP1BRESP(),  // out std_logic_vector(1 downto 0);
    .SAXIHP1BVALID(),  // out std_ulogic;
    .SAXIHP1RACOUNT(),  // out std_logic_vector(2 downto 0);
    .SAXIHP1RCOUNT(),  // out std_logic_vector(7 downto 0);
    .SAXIHP1RDATA(),  // out std_logic_vector(63 downto 0);
    .SAXIHP1RID(), 	 // out std_logic_vector(5 downto 0);
    .SAXIHP1RLAST(),  // out std_ulogic;
    .SAXIHP1RRESP(),  // out std_logic_vector(1 downto 0);
    .SAXIHP1RVALID(),  // out std_ulogic;
    .SAXIHP1WACOUNT(),  // out std_logic_vector(5 downto 0);
    .SAXIHP1WCOUNT(),  // out std_logic_vector(7 downto 0);
    .SAXIHP1WREADY(),  // out std_ulogic;
    .SAXIHP2ARESETN(),  // out std_ulogic;
    .SAXIHP2ARREADY(),  // out std_ulogic;
    .SAXIHP2AWREADY(),  // out std_ulogic;
    .SAXIHP2BID(), 	 // out std_logic_vector(5 downto 0);
    .SAXIHP2BRESP(),  // out std_logic_vector(1 downto 0);
    .SAXIHP2BVALID(),  // out std_ulogic;
    .SAXIHP2RACOUNT(),  // out std_logic_vector(2 downto 0);
    .SAXIHP2RCOUNT(),  // out std_logic_vector(7 downto 0);
    .SAXIHP2RDATA(),  // out std_logic_vector(63 downto 0);
    .SAXIHP2RID(), 	 // out std_logic_vector(5 downto 0);
    .SAXIHP2RLAST(),  // out std_ulogic;
    .SAXIHP2RRESP(),  // out std_logic_vector(1 downto 0);
    .SAXIHP2RVALID(),  // out std_ulogic;
    .SAXIHP2WACOUNT(),  // out std_logic_vector(5 downto 0);
    .SAXIHP2WCOUNT(),  // out std_logic_vector(7 downto 0);
    .SAXIHP2WREADY(),  // out std_ulogic;
    .SAXIHP3ARESETN(),  // out std_ulogic;
    .SAXIHP3ARREADY(),  // out std_ulogic;
    .SAXIHP3AWREADY(),  // out std_ulogic;
    .SAXIHP3BID(), 	 // out std_logic_vector(5 downto 0);
    .SAXIHP3BRESP(),  // out std_logic_vector(1 downto 0);
    .SAXIHP3BVALID(),  // out std_ulogic;
    .SAXIHP3RACOUNT(),  // out std_logic_vector(2 downto 0);
    .SAXIHP3RCOUNT(),  // out std_logic_vector(7 downto 0);
    .SAXIHP3RDATA(),  // out std_logic_vector(63 downto 0);
    .SAXIHP3RID(), 	 // out std_logic_vector(5 downto 0);
    .SAXIHP3RLAST(),  // out std_ulogic;
    .SAXIHP3RRESP(),  // out std_logic_vector(1 downto 0);
    .SAXIHP3RVALID(),  // out std_ulogic;
    .SAXIHP3WACOUNT(),  // out std_logic_vector(5 downto 0);
    .SAXIHP3WCOUNT(),  // out std_logic_vector(7 downto 0);
    .SAXIHP3WREADY(),  // out std_ulogic;
    .DDRA(DDR_Addr), 	// inout std_logic_vector(14 downto 0);
    .DDRBA(DDR_BankAddr), // inout std_logic_vector(2 downto 0);
    .DDRCASB(DDR_CAS_n), 	// inout std_ulogic;
    .DDRCKE(DDR_CKE), 	// inout std_ulogic;
    .DDRCKN(DDR_Clk_n), 	// inout std_ulogic;
    .DDRCKP(DDR_Clk), 	// inout std_ulogic;
    .DDRCSB(DDR_CS_n), 	// inout std_ulogic;
    .DDRDM(DDR_DM), 	// inout std_logic_vector(3 downto 0);
    .DDRDQ(DDR_DQ), 	// inout std_logic_vector(31 downto 0);
    .DDRDQSN(DDR_DQS_n), 	// inout std_logic_vector(3 downto 0);
    .DDRDQSP(DDR_DQS), 	// inout std_logic_vector(3 downto 0);
    .DDRDRSTB(DDR_DRSTB), 	// inout std_ulogic;
    .DDRODT(DDR_ODT), 	// inout std_ulogic;
    .DDRRASB(DDR_RAS_n), 	// inout std_ulogic;
    .DDRVRN(DDR_VRN), 	// inout std_ulogic;
    .DDRVRP(DDR_VRP), 	// inout std_ulogic;
    .DDRWEB(DDR_WEB), 	// inout std_ulogic;
    .MIO(MIO), 	// inout std_logic_vector(53 downto 0);
    .PSCLK(PS_CLK), 	// inout std_ulogic;
    .PSPORB(PS_PORB), 	// inout std_ulogic;
    .PSSRSTB(PS_SRSTB), 	// inout std_ulogic;
    .DDRARB(4'b0),	// in std_logic_vector(3 downto 0);
    .DMA0ACLK(1'b0), 		// in std_ulogic;
    .DMA0DAREADY(1'b0), 		// in std_ulogic;
    .DMA0DRLAST(1'b0), 		// in std_ulogic;
    .DMA0DRTYPE(2'b0),	// in std_logic_vector(1 downto 0);
    .DMA0DRVALID(1'b0), 		// in std_ulogic;
    .DMA1ACLK(1'b0), 		// in std_ulogic;
    .DMA1DAREADY(1'b0), 		// in std_ulogic;
    .DMA1DRLAST(1'b0), 		// in std_ulogic;
    .DMA1DRTYPE(2'b0),	// in std_logic_vector(1 downto 0);
    .DMA1DRVALID(1'b0), 		// in std_ulogic;
    .DMA2ACLK(1'b0), 		// in std_ulogic;
    .DMA2DAREADY(1'b0), 		// in std_ulogic;
    .DMA2DRLAST(1'b0), 		// in std_ulogic;
    .DMA2DRTYPE(2'b0),	// in std_logic_vector(1 downto 0);
    .DMA2DRVALID(1'b0), 		// in std_ulogic;
    .DMA3ACLK(1'b0), 		// in std_ulogic;
    .DMA3DAREADY(1'b0), 		// in std_ulogic;
    .DMA3DRLAST(1'b0), 		// in std_ulogic;
    .DMA3DRTYPE(2'b0),	// in std_logic_vector(1 downto 0);
    .DMA3DRVALID(1'b0), 		// in std_ulogic;
    .EMIOCAN0PHYRX(1'b0), 		// in std_ulogic;
    .EMIOCAN1PHYRX(1'b0), 		// in std_ulogic;
    .EMIOENET0EXTINTIN(1'b0), 		// in std_ulogic;
    .EMIOENET0GMIICOL(1'b0), 		// in std_ulogic;
    .EMIOENET0GMIICRS(1'b0), 		// in std_ulogic;
    .EMIOENET0GMIIRXCLK(1'b0), 		// in std_ulogic;
    .EMIOENET0GMIIRXD(8'b0),	// in std_logic_vector(7 downto 0);
    .EMIOENET0GMIIRXDV(1'b0), 		// in std_ulogic;
    .EMIOENET0GMIIRXER(1'b0), 		// in std_ulogic;
    .EMIOENET0GMIITXCLK(1'b0), 		// in std_ulogic;
    .EMIOENET0MDIOI(1'b0), 		// in std_ulogic;
    .EMIOENET1EXTINTIN(1'b0), 		// in std_ulogic;
    .EMIOENET1GMIICOL(1'b0), 		// in std_ulogic;
    .EMIOENET1GMIICRS(1'b0), 		// in std_ulogic;
    .EMIOENET1GMIIRXCLK(1'b0), 		// in std_ulogic;
    .EMIOENET1GMIIRXD(8'b0),	// in std_logic_vector(7 downto 0);
    .EMIOENET1GMIIRXDV(1'b0), 		// in std_ulogic;
    .EMIOENET1GMIIRXER(1'b0), 		// in std_ulogic;
    .EMIOENET1GMIITXCLK(1'b0), 		// in std_ulogic;
    .EMIOENET1MDIOI(1'b0), 		// in std_ulogic;
    .EMIOGPIOI(64'b0), 	// in std_logic_vector(63 downto 0);
    .EMIOI2C0SCLI(1'b0), 	// in std_ulogic;
    .EMIOI2C0SDAI(1'b0), 	// in std_ulogic;
    .EMIOI2C1SCLI(1'b0), 	// in std_ulogic;
    .EMIOI2C1SDAI(1'b0), 	// in std_ulogic;
    .EMIOPJTAGTCK(1'b0), 		// in std_ulogic;
    .EMIOPJTAGTDI(1'b0), 		// in std_ulogic;
    .EMIOPJTAGTMS(1'b0), 		// in std_ulogic;
    .EMIOSDIO0CDN(1'b0), 		// in std_ulogic;
    .EMIOSDIO0CLKFB(1'b0), 		// in std_ulogic;
    .EMIOSDIO0CMDI(1'b0), 		// in std_ulogic;
    .EMIOSDIO0DATAI(4'b0),	// in std_logic_vector(3 downto 0);
    .EMIOSDIO0WP(1'b0), 		// in std_ulogic;
    .EMIOSDIO1CDN(1'b0), 		// in std_ulogic;
    .EMIOSDIO1CLKFB(1'b0), 		// in std_ulogic;
    .EMIOSDIO1CMDI(1'b0), 		// in std_ulogic;
    .EMIOSDIO1DATAI(4'b0),	// in std_logic_vector(3 downto 0);
    .EMIOSDIO1WP(1'b0), 		// in std_ulogic;
    .EMIOSPI0MI(1'b0), 		// in std_ulogic;
    .EMIOSPI0SCLKI(1'b0), 		// in std_ulogic;
    .EMIOSPI0SI(1'b0), 		// in std_ulogic;
    .EMIOSPI0SSIN(1'b0), 		// in std_ulogic;
    .EMIOSPI1MI(1'b0), 		// in std_ulogic;
    .EMIOSPI1SCLKI(1'b0), 		// in std_ulogic;
    .EMIOSPI1SI(1'b0), 		// in std_ulogic;
    .EMIOSPI1SSIN(1'b0), 		// in std_ulogic;
    .EMIOSRAMINTIN(1'b0), 		// in std_ulogic;
    .EMIOTRACECLK(1'b0), 		// in std_ulogic;
    .EMIOTTC0CLKI(3'b0),	// in std_logic_vector(2 downto 0);
    .EMIOTTC1CLKI(3'b0),	// in std_logic_vector(2 downto 0);
    .EMIOUART0CTSN(1'b0), 		// in std_ulogic;
    .EMIOUART0DCDN(1'b0), 		// in std_ulogic;
    .EMIOUART0DSRN(1'b0), 		// in std_ulogic;
    .EMIOUART0RIN(1'b0), 		// in std_ulogic;
    .EMIOUART0RX(1'b0), 		// in std_ulogic;
    .EMIOUART1CTSN(1'b0), 		// in std_ulogic;
    .EMIOUART1DCDN(1'b0), 		// in std_ulogic;
    .EMIOUART1DSRN(1'b0), 		// in std_ulogic;
    .EMIOUART1RIN(1'b0), 		// in std_ulogic;
    .EMIOUART1RX(1'b0), 		// in std_ulogic;
    .EMIOUSB0VBUSPWRFAULT(1'b0), 		// in std_ulogic;
    .EMIOUSB1VBUSPWRFAULT(1'b0), 		// in std_ulogic;
    .EMIOWDTCLKI(1'b0), 		// in std_ulogic;
    .EVENTEVENTI(1'b0), 		// in std_ulogic;
    .FCLKCLKTRIGN(4'b0),	// in std_logic_vector(3 downto 0);
    .FPGAIDLEN(1'b0), 		// in std_ulogic;
    .FTMDTRACEINATID(4'b0),	// in std_logic_vector(3 downto 0);
    .FTMDTRACEINCLOCK(1'b0), 		// in std_ulogic;
    .FTMDTRACEINDATA(32'b0),	// in std_logic_vector(31 downto 0);
    .FTMDTRACEINVALID(1'b0), 		// in std_ulogic;
    .FTMTF2PDEBUG(32'b0),	// in std_logic_vector(31 downto 0);
    .FTMTF2PTRIG(4'b0),	// in std_logic_vector(3 downto 0);
    .FTMTP2FTRIGACK(4'b0),	// in std_logic_vector(3 downto 0);
    .IRQF2P({19'b0,CONFIG_IRQ}),	// in std_logic_vector(19 downto 0);
    .MAXIGP1ACLK(1'b0), 	// in std_ulogic;
    .MAXIGP1ARREADY(1'b0), // in std_ulogic;
    .MAXIGP1AWREADY(1'b0), // in std_ulogic;
    .MAXIGP1BID(12'b0), 	// in std_logic_vector(11 downto 0);
    .MAXIGP1BRESP(2'b0), // in std_logic_vector(1 downto 0);
    .MAXIGP1BVALID(1'b0), // in std_ulogic;
    .MAXIGP1RDATA(32'b0), // in std_logic_vector(31 downto 0);
    .MAXIGP1RID(12'b0), 	// in std_logic_vector(11 downto 0);
    .MAXIGP1RLAST(1'b0), // in std_ulogic;
    .MAXIGP1RRESP(2'b0), // in std_logic_vector(1 downto 0);
    .MAXIGP1RVALID(1'b0), // in std_ulogic;
    .MAXIGP1WREADY(1'b0), // in std_ulogic;
    .SAXIGP0ACLK(1'b0), 		// in std_ulogic;
    .SAXIGP0ARADDR(32'b0),	// in std_logic_vector(31 downto 0);
    .SAXIGP0ARBURST(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP0ARCACHE(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP0ARID(6'b0),	// in std_logic_vector(5 downto 0);
    .SAXIGP0ARLEN(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP0ARLOCK(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP0ARPROT(3'b0),	// in std_logic_vector(2 downto 0);
    .SAXIGP0ARQOS(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP0ARSIZE(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP0ARVALID(1'b0), 		// in std_ulogic;
    .SAXIGP0AWADDR(32'b0),	// in std_logic_vector(31 downto 0);
    .SAXIGP0AWBURST(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP0AWCACHE(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP0AWID(6'b0),	// in std_logic_vector(5 downto 0);
    .SAXIGP0AWLEN(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP0AWLOCK(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP0AWPROT(3'b0),	// in std_logic_vector(2 downto 0);
    .SAXIGP0AWQOS(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP0AWSIZE(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP0AWVALID(1'b0), 		// in std_ulogic;
    .SAXIGP0BREADY(1'b0), 		// in std_ulogic;
    .SAXIGP0RREADY(1'b0), 		// in std_ulogic;
    .SAXIGP0WDATA(32'b0),	// in std_logic_vector(31 downto 0);
    .SAXIGP0WID(6'b0),	// in std_logic_vector(5 downto 0);
    .SAXIGP0WLAST(1'b0), 		// in std_ulogic;
    .SAXIGP0WSTRB(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP0WVALID(1'b0), 		// in std_ulogic;
    .SAXIGP1ACLK(1'b0), 		// in std_ulogic;
    .SAXIGP1ARADDR(32'b0),	// in std_logic_vector(31 downto 0);
    .SAXIGP1ARBURST(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP1ARCACHE(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP1ARID(6'b0),	// in std_logic_vector(5 downto 0);
    .SAXIGP1ARLEN(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP1ARLOCK(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP1ARPROT(3'b0),	// in std_logic_vector(2 downto 0);
    .SAXIGP1ARQOS(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP1ARSIZE(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP1ARVALID(1'b0), 		// in std_ulogic;
    .SAXIGP1AWADDR(32'b0),	// in std_logic_vector(31 downto 0);
    .SAXIGP1AWBURST(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP1AWCACHE(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP1AWID(6'b0),	// in std_logic_vector(5 downto 0);
    .SAXIGP1AWLEN(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP1AWLOCK(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP1AWPROT(3'b0),	// in std_logic_vector(2 downto 0);
    .SAXIGP1AWQOS(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP1AWSIZE(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP1AWVALID(1'b0), 		// in std_ulogic;
    .SAXIGP1BREADY(1'b0), 		// in std_ulogic;
    .SAXIGP1RREADY(1'b0), 		// in std_ulogic;
    .SAXIGP1WDATA(32'b0),	// in std_logic_vector(31 downto 0);
    .SAXIGP1WID(6'b0),	// in std_logic_vector(5 downto 0);
    .SAXIGP1WLAST(1'b0), 		// in std_ulogic;
    .SAXIGP1WSTRB(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP1WVALID(1'b0), 		// in std_ulogic;
    .SAXIHP1ACLK(1'b0), 	// in std_ulogic;
    .SAXIHP1ARADDR(32'b0), // in std_logic_vector(31 downto 0);
    .SAXIHP1ARBURST(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP1ARCACHE(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP1ARID(6'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIHP1ARLEN(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP1ARLOCK(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP1ARPROT(3'b0), // in std_logic_vector(2 downto 0);
    .SAXIHP1ARQOS(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP1ARSIZE(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP1ARVALID(1'b0), // in std_ulogic;
    .SAXIHP1AWADDR(32'b0), // in std_logic_vector(31 downto 0);
    .SAXIHP1AWBURST(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP1AWCACHE(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP1AWID(6'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIHP1AWLEN(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP1AWLOCK(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP1AWPROT(3'b0), // in std_logic_vector(2 downto 0);
    .SAXIHP1AWQOS(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP1AWSIZE(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP1AWVALID(1'b0), // in std_ulogic;
    .SAXIHP1BREADY(1'b0), // in std_ulogic;
    .SAXIHP1RDISSUECAP1EN(1'b0), 		// in std_ulogic;
    .SAXIHP1RREADY(1'b0), // in std_ulogic;
    .SAXIHP1WDATA(64'b0), // in std_logic_vector(63 downto 0);
    .SAXIHP1WID(6'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIHP1WLAST(1'b0), // in std_ulogic;
    .SAXIHP1WRISSUECAP1EN(1'b0), 		// in std_ulogic;
    .SAXIHP1WSTRB(8'b0), // in std_logic_vector(7 downto 0);
    .SAXIHP1WVALID(1'b0), // in std_ulogic;
    .SAXIHP2ACLK(1'b0), 	// in std_ulogic;
    .SAXIHP2ARADDR(32'b0), // in std_logic_vector(31 downto 0);
    .SAXIHP2ARBURST(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP2ARCACHE(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP2ARID(6'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIHP2ARLEN(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP2ARLOCK(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP2ARPROT(3'b0), // in std_logic_vector(2 downto 0);
    .SAXIHP2ARQOS(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP2ARSIZE(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP2ARVALID(1'b0), // in std_ulogic;
    .SAXIHP2AWADDR(32'b0), // in std_logic_vector(31 downto 0);
    .SAXIHP2AWBURST(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP2AWCACHE(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP2AWID(6'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIHP2AWLEN(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP2AWLOCK(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP2AWPROT(3'b0), // in std_logic_vector(2 downto 0);
    .SAXIHP2AWQOS(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP2AWSIZE(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP2AWVALID(1'b0), // in std_ulogic;
    .SAXIHP2BREADY(1'b0), // in std_ulogic;
    .SAXIHP2RDISSUECAP1EN(1'b0), 		// in std_ulogic;
    .SAXIHP2RREADY(1'b0), // in std_ulogic;
    .SAXIHP2WDATA(64'b0), // in std_logic_vector(63 downto 0);
    .SAXIHP2WID(6'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIHP2WLAST(1'b0), // in std_ulogic;
    .SAXIHP2WRISSUECAP1EN(1'b0), 		// in std_ulogic;
    .SAXIHP2WSTRB(8'b0), // in std_logic_vector(7 downto 0);
    .SAXIHP2WVALID(1'b0), // in std_ulogic;
    .SAXIHP3ACLK(1'b0), 	// in std_ulogic;
    .SAXIHP3ARADDR(32'b0), // in std_logic_vector(31 downto 0);
    .SAXIHP3ARBURST(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP3ARCACHE(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP3ARID(6'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIHP3ARLEN(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP3ARLOCK(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP3ARPROT(3'b0), // in std_logic_vector(2 downto 0);
    .SAXIHP3ARQOS(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP3ARSIZE(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP3ARVALID(1'b0), // in std_ulogic;
    .SAXIHP3AWADDR(32'b0), // in std_logic_vector(31 downto 0);
    .SAXIHP3AWBURST(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP3AWCACHE(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP3AWID(6'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIHP3AWLEN(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP3AWLOCK(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP3AWPROT(3'b0), // in std_logic_vector(2 downto 0);
    .SAXIHP3AWQOS(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP3AWSIZE(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP3AWVALID(1'b0), // in std_ulogic;
    .SAXIHP3BREADY(1'b0), // in std_ulogic;
    .SAXIHP3RDISSUECAP1EN(1'b0), 		// in std_ulogic;
    .SAXIHP3RREADY(1'b0), // in std_ulogic;
    .SAXIHP3WDATA(64'b0), // in std_logic_vector(63 downto 0);
    .SAXIHP3WID(6'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIHP3WLAST(1'b0), // in std_ulogic;
    .SAXIHP3WRISSUECAP1EN(1'b0), 		// in std_ulogic;
    .SAXIHP3WSTRB(8'b0), // in std_logic_vector(7 downto 0);
    .SAXIHP3WVALID(1'b0)	// in std_ulogic;
  );
endmodule
