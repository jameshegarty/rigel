module incif_1uint32_CEtable__0x45fd16f0(input CLK, input CE, input [32:0] process_input, output [31:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [31:0] unnamedcast36583USEDMULTIPLEcast;assign unnamedcast36583USEDMULTIPLEcast = (process_input[31:0]); 
  assign process_output = (((process_input[32]))?({(unnamedcast36583USEDMULTIPLEcast+(32'd1))}):(unnamedcast36583USEDMULTIPLEcast));
  // function: process pure=true delay=0
endmodule

module RegBy_incif_1uint32_CEtable__0x45fd16f0_CEtrue_initnil(input CLK, input set_valid, input CE, input [31:0] set_inp, input setby_valid, input setby_inp, output [31:0] SETBY_OUTPUT, output [31:0] GET_OUTPUT);
parameter INSTANCE_NAME="INST";
  reg [31:0] R;
  wire [31:0] regby_inner_process_output;
  always @(posedge CLK) begin if(set_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(setby_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,set_valid})+({4'b0,setby_valid})) > 5'd1) begin $display("error, function 'set' on instance 'R' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [32:0] unnamedcallArbitrate36615USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate36615USEDMULTIPLEcallArbitrate = {(set_valid||setby_valid),((set_valid)?(set_inp):(regby_inner_process_output))}; 
    always @ (posedge CLK) begin if ((unnamedcallArbitrate36615USEDMULTIPLEcallArbitrate[32]) && CE) begin R <= (unnamedcallArbitrate36615USEDMULTIPLEcallArbitrate[31:0]); end end
  assign SETBY_OUTPUT = regby_inner_process_output;
  assign GET_OUTPUT = R;
  // function: set pure=false ONLY WIRE
  // function: setby pure=false ONLY WIRE
  // function: get pure=true ONLY WIRE
  incif_1uint32_CEtable__0x45fd16f0 #(.INSTANCE_NAME({INSTANCE_NAME,"_regby_inner"})) regby_inner(.CLK(CLK), .CE(CE), .process_input({setby_inp,R}), .process_output(regby_inner_process_output));
endmodule

module Underflow_Auint8_2_1__4_1__count76800_cycles6087906_toosoonnil_UStrue(input CLK, input ready_downstream, output ready, input reset, input [64:0] process_input, output [64:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire [31:0] cycleCount_GET_OUTPUT;
  wire unnamedbinop37596USEDMULTIPLEbinop;assign unnamedbinop37596USEDMULTIPLEbinop = {((cycleCount_GET_OUTPUT)>((32'd6087906)))}; 
  assign ready = {(ready_downstream||unnamedbinop37596USEDMULTIPLEbinop)};
  wire unnamedbinop37598USEDMULTIPLEbinop;assign unnamedbinop37598USEDMULTIPLEbinop = {({(ready_downstream||reset)}||unnamedbinop37596USEDMULTIPLEbinop)}; 
  wire [31:0] outputCount_GET_OUTPUT;
  wire unnamedcast37590USEDMULTIPLEcast;assign unnamedcast37590USEDMULTIPLEcast = (process_input[64]); 
  wire unnamedunary37618USEDMULTIPLEunary;assign unnamedunary37618USEDMULTIPLEunary = {(~reset)}; 
  wire [31:0] outputCount_SETBY_OUTPUT;
  wire [31:0] cycleCount_SETBY_OUTPUT;
  assign process_output = {{({({(unnamedbinop37596USEDMULTIPLEbinop&&{((outputCount_GET_OUTPUT)<((32'd76800)))})}||{({(~unnamedbinop37596USEDMULTIPLEbinop)}&&unnamedcast37590USEDMULTIPLEcast)})}&&unnamedunary37618USEDMULTIPLEunary)},((unnamedbinop37596USEDMULTIPLEbinop)?((64'd3735928559)):((process_input[63:0])))};
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  RegBy_incif_1uint32_CEtable__0x45fd16f0_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_outputCount"})) outputCount(.CLK(CLK), .set_valid(reset), .CE(unnamedbinop37598USEDMULTIPLEbinop), .set_inp((32'd0)), .setby_valid(unnamedunary37618USEDMULTIPLEunary), .setby_inp({(ready_downstream&&{(unnamedcast37590USEDMULTIPLEcast||unnamedbinop37596USEDMULTIPLEbinop)})}), .SETBY_OUTPUT(outputCount_SETBY_OUTPUT), .GET_OUTPUT(outputCount_GET_OUTPUT));
  RegBy_incif_1uint32_CEtable__0x45fd16f0_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_cycleCount"})) cycleCount(.CLK(CLK), .set_valid(reset), .CE((1'd1)), .set_inp((32'd0)), .setby_valid(unnamedunary37618USEDMULTIPLEunary), .setby_inp((1'd1)), .SETBY_OUTPUT(cycleCount_SETBY_OUTPUT), .GET_OUTPUT(cycleCount_GET_OUTPUT));
endmodule

module incif_wrapuint8_127_incnil(input CLK, input CE, input [8:0] process_input, output [7:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [7:0] unnamedcast693USEDMULTIPLEcast;assign unnamedcast693USEDMULTIPLEcast = (process_input[7:0]); 
  assign process_output = (((process_input[8]))?((({(unnamedcast693USEDMULTIPLEcast==(8'd127))})?((8'd0)):({(unnamedcast693USEDMULTIPLEcast+(8'd1))}))):(unnamedcast693USEDMULTIPLEcast));
  // function: process pure=true delay=0
endmodule

module RegBy_incif_wrapuint8_127_incnil_CEtrue_initnil(input CLK, input set_valid, input CE, input [7:0] set_inp, input setby_valid, input setby_inp, output [7:0] SETBY_OUTPUT, output [7:0] GET_OUTPUT);
parameter INSTANCE_NAME="INST";
  reg [7:0] R;
  wire [7:0] regby_inner_process_output;
  always @(posedge CLK) begin if(set_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(setby_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,set_valid})+({4'b0,setby_valid})) > 5'd1) begin $display("error, function 'set' on instance 'R' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [8:0] unnamedcallArbitrate744USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate744USEDMULTIPLEcallArbitrate = {(set_valid||setby_valid),((set_valid)?(set_inp):(regby_inner_process_output))}; 
    always @ (posedge CLK) begin if ((unnamedcallArbitrate744USEDMULTIPLEcallArbitrate[8]) && CE) begin R <= (unnamedcallArbitrate744USEDMULTIPLEcallArbitrate[7:0]); end end
  assign SETBY_OUTPUT = regby_inner_process_output;
  assign GET_OUTPUT = R;
  // function: set pure=false ONLY WIRE
  // function: setby pure=false ONLY WIRE
  // function: get pure=true ONLY WIRE
  incif_wrapuint8_127_incnil #(.INSTANCE_NAME({INSTANCE_NAME,"_regby_inner"})) regby_inner(.CLK(CLK), .CE(CE), .process_input({setby_inp,R}), .process_output(regby_inner_process_output));
endmodule

module fifo_uint8_128(input CLK, input popFront_valid, input CE_pop, output [7:0] popFront, output [7:0] size, input pushBackReset_valid, input CE_push, output ready, input pushBack_valid, input [7:0] pushBack_input, input popFrontReset_valid, output hasData);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(popFront_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'popFront'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(pushBackReset_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'pushBackReset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(pushBack_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'pushBack'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(popFrontReset_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'popFrontReset'", INSTANCE_NAME);  end end
  wire [7:0] readAddr_GET_OUTPUT;
  wire [6:0] unnamedcast820USEDMULTIPLEcast;assign unnamedcast820USEDMULTIPLEcast = readAddr_GET_OUTPUT[6:0]; 
  wire fifo1_READ_OUTPUT;
  wire fifo2_READ_OUTPUT;
  wire fifo3_READ_OUTPUT;
  wire fifo4_READ_OUTPUT;
  wire fifo5_READ_OUTPUT;
  wire fifo6_READ_OUTPUT;
  wire fifo7_READ_OUTPUT;
  wire fifo8_READ_OUTPUT;
  wire [7:0] writeAddr_GET_OUTPUT;
  wire unnamedunary767USEDMULTIPLEunary;assign unnamedunary767USEDMULTIPLEunary = {(~{(writeAddr_GET_OUTPUT==readAddr_GET_OUTPUT)})}; 
  always @(posedge CLK) begin if(unnamedunary767USEDMULTIPLEunary == 1'b0 && popFront_valid==1'b1 && CE_pop==1'b1) begin $display("%s: attempting to pop from an empty fifo",INSTANCE_NAME);$finish();  end end
  wire [7:0] readAddr_SETBY_OUTPUT;
  assign popFront = {fifo8_READ_OUTPUT,fifo7_READ_OUTPUT,fifo6_READ_OUTPUT,fifo5_READ_OUTPUT,fifo4_READ_OUTPUT,fifo3_READ_OUTPUT,fifo2_READ_OUTPUT,fifo1_READ_OUTPUT};
  wire [7:0] unnamedselect758USEDMULTIPLEselect;assign unnamedselect758USEDMULTIPLEselect = (({((writeAddr_GET_OUTPUT)<(readAddr_GET_OUTPUT))})?({({((8'd128)-readAddr_GET_OUTPUT)}+writeAddr_GET_OUTPUT)}):({(writeAddr_GET_OUTPUT-readAddr_GET_OUTPUT)})); 
  assign size = unnamedselect758USEDMULTIPLEselect;
  reg readyReg;
    always @ (posedge CLK) begin readyReg <= {((unnamedselect758USEDMULTIPLEselect)<((8'd125)))}; end
  assign ready = readyReg;
  always @(posedge CLK) begin if({((unnamedselect758USEDMULTIPLEselect)<((8'd126)))} == 1'b0 && pushBack_valid==1'b1 && CE_push==1'b1) begin $display("%s: attempting to push to a full fifo",INSTANCE_NAME);$finish();  end end
  wire [7:0] writeAddr_SETBY_OUTPUT;
  wire [6:0] unnamedcast775USEDMULTIPLEcast;assign unnamedcast775USEDMULTIPLEcast = writeAddr_GET_OUTPUT[6:0]; 
  assign hasData = unnamedunary767USEDMULTIPLEunary;
  // function: popFront pure=false delay=0
  // function: size pure=true delay=0
  // function: pushBackReset pure=false delay=0
  // function: ready pure=true delay=0
  // function: pushBack pure=false delay=0
  // function: popFrontReset pure=false delay=0
  // function: hasData pure=true delay=0
  RegBy_incif_wrapuint8_127_incnil_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_writeAddr"})) writeAddr(.CLK(CLK), .set_valid(pushBackReset_valid), .CE(CE_push), .set_inp((8'd0)), .setby_valid(pushBack_valid), .setby_inp((1'd1)), .SETBY_OUTPUT(writeAddr_SETBY_OUTPUT), .GET_OUTPUT(writeAddr_GET_OUTPUT));
  RegBy_incif_wrapuint8_127_incnil_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_readAddr"})) readAddr(.CLK(CLK), .set_valid(popFrontReset_valid), .CE(CE_pop), .set_inp((8'd0)), .setby_valid(popFront_valid), .setby_inp((1'd1)), .SETBY_OUTPUT(readAddr_SETBY_OUTPUT), .GET_OUTPUT(readAddr_GET_OUTPUT));
  wire [7:0] fifo1_writeInput = {pushBack_input[0:0],unnamedcast775USEDMULTIPLEcast};
wire fifo1_writeOut;
RAM128X1D fifo1  (
  .WCLK(CLK),
  .D(fifo1_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo1_writeOut),
  .DPO(fifo1_READ_OUTPUT),
  .A(fifo1_writeInput[6:0]),
  .DPRA(unnamedcast820USEDMULTIPLEcast));

  wire [7:0] fifo2_writeInput = {pushBack_input[1:1],unnamedcast775USEDMULTIPLEcast};
wire fifo2_writeOut;
RAM128X1D fifo2  (
  .WCLK(CLK),
  .D(fifo2_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo2_writeOut),
  .DPO(fifo2_READ_OUTPUT),
  .A(fifo2_writeInput[6:0]),
  .DPRA(unnamedcast820USEDMULTIPLEcast));

  wire [7:0] fifo3_writeInput = {pushBack_input[2:2],unnamedcast775USEDMULTIPLEcast};
wire fifo3_writeOut;
RAM128X1D fifo3  (
  .WCLK(CLK),
  .D(fifo3_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo3_writeOut),
  .DPO(fifo3_READ_OUTPUT),
  .A(fifo3_writeInput[6:0]),
  .DPRA(unnamedcast820USEDMULTIPLEcast));

  wire [7:0] fifo4_writeInput = {pushBack_input[3:3],unnamedcast775USEDMULTIPLEcast};
wire fifo4_writeOut;
RAM128X1D fifo4  (
  .WCLK(CLK),
  .D(fifo4_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo4_writeOut),
  .DPO(fifo4_READ_OUTPUT),
  .A(fifo4_writeInput[6:0]),
  .DPRA(unnamedcast820USEDMULTIPLEcast));

  wire [7:0] fifo5_writeInput = {pushBack_input[4:4],unnamedcast775USEDMULTIPLEcast};
wire fifo5_writeOut;
RAM128X1D fifo5  (
  .WCLK(CLK),
  .D(fifo5_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo5_writeOut),
  .DPO(fifo5_READ_OUTPUT),
  .A(fifo5_writeInput[6:0]),
  .DPRA(unnamedcast820USEDMULTIPLEcast));

  wire [7:0] fifo6_writeInput = {pushBack_input[5:5],unnamedcast775USEDMULTIPLEcast};
wire fifo6_writeOut;
RAM128X1D fifo6  (
  .WCLK(CLK),
  .D(fifo6_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo6_writeOut),
  .DPO(fifo6_READ_OUTPUT),
  .A(fifo6_writeInput[6:0]),
  .DPRA(unnamedcast820USEDMULTIPLEcast));

  wire [7:0] fifo7_writeInput = {pushBack_input[6:6],unnamedcast775USEDMULTIPLEcast};
wire fifo7_writeOut;
RAM128X1D fifo7  (
  .WCLK(CLK),
  .D(fifo7_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo7_writeOut),
  .DPO(fifo7_READ_OUTPUT),
  .A(fifo7_writeInput[6:0]),
  .DPRA(unnamedcast820USEDMULTIPLEcast));

  wire [7:0] fifo8_writeInput = {pushBack_input[7:7],unnamedcast775USEDMULTIPLEcast};
wire fifo8_writeOut;
RAM128X1D fifo8  (
  .WCLK(CLK),
  .D(fifo8_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo8_writeOut),
  .DPO(fifo8_READ_OUTPUT),
  .A(fifo8_writeInput[6:0]),
  .DPRA(unnamedcast820USEDMULTIPLEcast));

endmodule

module fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128(input CLK, input load_valid, input load_CE, output [8:0] load_output, input store_reset_valid, input store_CE, output store_ready, input load_reset_valid, input store_valid, input [7:0] store_input);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(load_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_reset_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(load_reset_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store'", INSTANCE_NAME);  end end
  wire FIFO_hasData;
  wire [7:0] FIFO_popFront;
  assign load_output = {FIFO_hasData,FIFO_popFront};
  wire FIFO_ready;
  assign store_ready = FIFO_ready;
  // function: load pure=false delay=0
  // function: store_reset pure=false delay=0
  // function: store_ready pure=true delay=0
  // function: load_reset pure=false delay=0
  // function: store pure=false delay=0
  fifo_uint8_128 #(.INSTANCE_NAME({INSTANCE_NAME,"_FIFO"})) FIFO(.CLK(CLK), .popFront_valid({(FIFO_hasData&&load_valid)}), .CE_pop(load_CE), .popFront(FIFO_popFront), .size(FIFO_size), .pushBackReset_valid(store_reset_valid), .CE_push(store_CE), .ready(FIFO_ready), .pushBack_valid(store_valid), .pushBack_input(store_input), .popFrontReset_valid(load_reset_valid), .hasData(FIFO_hasData));
endmodule

module LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128(input CLK, input load_valid, input load_CE, input load_input, output [8:0] load_output, input store_reset_valid, input store_CE, output store_ready, output load_ready, input load_reset, input store_valid, input [7:0] store_input);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(load_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_reset_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(load_reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store'", INSTANCE_NAME);  end end
  wire unnamedcast1079USEDMULTIPLEcast;assign unnamedcast1079USEDMULTIPLEcast = load_input; 
  wire [8:0] LiftDecimate_load_output;
  reg [7:0] unnamedcast1082_delay1_validunnamednull0_CEload_CE;  always @ (posedge CLK) begin if (load_CE) begin unnamedcast1082_delay1_validunnamednull0_CEload_CE <= (LiftDecimate_load_output[7:0]); end end
  reg unnamedbinop1087_delay1_validunnamednull0_CEload_CE;  always @ (posedge CLK) begin if (load_CE) begin unnamedbinop1087_delay1_validunnamednull0_CEload_CE <= {((LiftDecimate_load_output[8])&&unnamedcast1079USEDMULTIPLEcast)}; end end
  assign load_output = {unnamedbinop1087_delay1_validunnamednull0_CEload_CE,unnamedcast1082_delay1_validunnamednull0_CEload_CE};
  wire LiftDecimate_store_ready;
  assign store_ready = LiftDecimate_store_ready;
  assign load_ready = (1'd1);
  // function: load pure=false delay=1
  // function: store_reset pure=false delay=0
  // function: store_ready pure=true delay=0
  // function: load_ready pure=true delay=0
  // function: load_reset pure=false delay=0
  // function: store pure=false delay=0
  fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128 #(.INSTANCE_NAME({INSTANCE_NAME,"_LiftDecimate"})) LiftDecimate(.CLK(CLK), .load_valid({(unnamedcast1079USEDMULTIPLEcast&&load_valid)}), .load_CE(load_CE), .load_output(LiftDecimate_load_output), .store_reset_valid(store_reset_valid), .store_CE(store_CE), .store_ready(LiftDecimate_store_ready), .load_reset_valid(load_reset), .store_valid(store_valid), .store_input(store_input));
endmodule

module RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128(input CLK, input load_valid, input load_CE, input load_input, output [8:0] load_output, input store_reset, input CE, output store_ready, output load_ready, input load_reset, input store_valid, input [8:0] store_input, output store_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(load_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(load_reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store'", INSTANCE_NAME);  end end
  wire [8:0] RunIffReady_load_output;
  assign load_output = RunIffReady_load_output;
  wire RunIffReady_store_ready;
  assign store_ready = RunIffReady_store_ready;
  wire RunIffReady_load_ready;
  assign load_ready = RunIffReady_load_ready;
  wire unnamedbinop1158USEDMULTIPLEbinop;assign unnamedbinop1158USEDMULTIPLEbinop = {({(RunIffReady_store_ready&&(store_input[8]))}&&store_valid)}; 
  assign store_output = {unnamedbinop1158USEDMULTIPLEbinop};
  // function: load pure=false delay=1
  // function: store_reset pure=false delay=0
  // function: store_ready pure=true delay=0
  // function: load_ready pure=true delay=0
  // function: load_reset pure=false delay=0
  // function: store pure=false delay=0
  LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128 #(.INSTANCE_NAME({INSTANCE_NAME,"_RunIffReady"})) RunIffReady(.CLK(CLK), .load_valid(load_valid), .load_CE(load_CE), .load_input(load_input), .load_output(RunIffReady_load_output), .store_reset_valid(store_reset), .store_CE(CE), .store_ready(RunIffReady_store_ready), .load_ready(RunIffReady_load_ready), .load_reset(load_reset), .store_valid(unnamedbinop1158USEDMULTIPLEbinop), .store_input((store_input[7:0])));
endmodule

module ShiftRegister_1_CEtrue_TY1(input CLK, input pushPop_valid, input CE, input sr_input, output pushPop_out, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'pushPop'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  reg SR1;
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR1' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR1' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR1' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate276USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate276USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(sr_input):((1'd0)))}; 
    always @ (posedge CLK) begin if ((unnamedcallArbitrate276USEDMULTIPLEcallArbitrate[1]) && CE) begin SR1 <= (unnamedcallArbitrate276USEDMULTIPLEcallArbitrate[0]); end end
  assign pushPop_out = SR1;
  // function: pushPop pure=false delay=0
  // function: reset pure=false delay=0
endmodule

module ShiftRegister_0_CEtrue_TY1(input CLK, input CE, input sr_input, output pushPop_out);
parameter INSTANCE_NAME="INST";
  assign pushPop_out = sr_input;
  // function: pushPop pure=true delay=0
  // function: reset pure=true delay=0
endmodule

module LiftHandshake_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128(input CLK, input load_input, output [8:0] load_output, input store_reset, input store_ready_downstream, output store_ready, input load_ready_downstream, output load_ready, input load_reset, input [8:0] store_input, output store_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire unnamedunary1195USEDMULTIPLEunary;assign unnamedunary1195USEDMULTIPLEunary = {(~load_reset)}; 
  wire unnamedbinop1194USEDMULTIPLEbinop;assign unnamedbinop1194USEDMULTIPLEbinop = {(load_reset||load_ready_downstream)}; 
  wire [8:0] inner_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128_load_output;
  wire load_validBitDelay_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128_pushPop_out;
  wire [8:0] unnamedtuple1205USEDMULTIPLEtuple;assign unnamedtuple1205USEDMULTIPLEtuple = {{((inner_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128_load_output[8])&&load_validBitDelay_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128_pushPop_out)},(inner_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128_load_output[7:0])}; 
  always @(posedge CLK) begin if({(~{((unnamedtuple1205USEDMULTIPLEtuple[8])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: output valid bit should not be X!",INSTANCE_NAME); end end
  always @(posedge CLK) begin if({(~{(load_input===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign load_output = unnamedtuple1205USEDMULTIPLEtuple;
  wire unnamedbinop1223USEDMULTIPLEbinop;assign unnamedbinop1223USEDMULTIPLEbinop = {(store_reset||store_ready_downstream)}; 
  wire inner_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128_store_ready;
  assign store_ready = {(inner_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128_store_ready&&store_ready_downstream)};
  wire inner_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128_load_ready;
  assign load_ready = {(inner_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128_load_ready&&load_ready_downstream)};
  wire unnamedunary1224USEDMULTIPLEunary;assign unnamedunary1224USEDMULTIPLEunary = {(~store_reset)}; 
  wire [0:0] inner_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128_store_output;
  wire store_validBitDelay_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128_pushPop_out;
  wire [0:0] unnamedtuple1234USEDMULTIPLEtuple;assign unnamedtuple1234USEDMULTIPLEtuple = {{(inner_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128_store_output&&store_validBitDelay_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128_pushPop_out)}}; 
  always @(posedge CLK) begin if({(~{(unnamedtuple1234USEDMULTIPLEtuple===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: output valid bit should not be X!",INSTANCE_NAME); end end
  always @(posedge CLK) begin if({(~{((store_input[8])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign store_output = unnamedtuple1234USEDMULTIPLEtuple;
  // function: load pure=false ONLY WIRE
  // function: store_reset pure=false ONLY WIRE
  // function: store_ready pure=true ONLY WIRE
  // function: load_ready pure=true ONLY WIRE
  // function: load_reset pure=false ONLY WIRE
  // function: store pure=false ONLY WIRE
  RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128 #(.INSTANCE_NAME({INSTANCE_NAME,"_inner_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128"})) inner_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128(.CLK(CLK), .load_valid(unnamedunary1195USEDMULTIPLEunary), .load_CE(unnamedbinop1194USEDMULTIPLEbinop), .load_input(load_input), .load_output(inner_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128_load_output), .store_reset(store_reset), .CE(unnamedbinop1223USEDMULTIPLEbinop), .store_ready(inner_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128_store_ready), .load_ready(inner_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128_load_ready), .load_reset(load_reset), .store_valid(unnamedunary1224USEDMULTIPLEunary), .store_input(store_input), .store_output(inner_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128_store_output));
  ShiftRegister_1_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_load_validBitDelay_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128"})) load_validBitDelay_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128(.CLK(CLK), .pushPop_valid(unnamedunary1195USEDMULTIPLEunary), .CE(unnamedbinop1194USEDMULTIPLEbinop), .sr_input((1'd1)), .pushPop_out(load_validBitDelay_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128_pushPop_out), .reset(load_reset));
  ShiftRegister_0_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_store_validBitDelay_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128"})) store_validBitDelay_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128(.CLK(CLK), .CE(unnamedbinop1223USEDMULTIPLEbinop), .sr_input((1'd1)), .pushPop_out(store_validBitDelay_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128_pushPop_out));
endmodule

module fifo__uint8_uint16__128(input CLK, input popFront_valid, input CE_pop, output [23:0] popFront, output [7:0] size, input pushBackReset_valid, input CE_push, output ready, input pushBack_valid, input [23:0] pushBack_input, input popFrontReset_valid, output hasData);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(popFront_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'popFront'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(pushBackReset_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'pushBackReset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(pushBack_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'pushBack'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(popFrontReset_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'popFrontReset'", INSTANCE_NAME);  end end
  wire [7:0] readAddr_GET_OUTPUT;
  wire [6:0] unnamedcast35117USEDMULTIPLEcast;assign unnamedcast35117USEDMULTIPLEcast = readAddr_GET_OUTPUT[6:0]; 
  wire fifo1_READ_OUTPUT;
  wire fifo2_READ_OUTPUT;
  wire fifo3_READ_OUTPUT;
  wire fifo4_READ_OUTPUT;
  wire fifo5_READ_OUTPUT;
  wire fifo6_READ_OUTPUT;
  wire fifo7_READ_OUTPUT;
  wire fifo8_READ_OUTPUT;
  wire fifo9_READ_OUTPUT;
  wire fifo10_READ_OUTPUT;
  wire fifo11_READ_OUTPUT;
  wire fifo12_READ_OUTPUT;
  wire fifo13_READ_OUTPUT;
  wire fifo14_READ_OUTPUT;
  wire fifo15_READ_OUTPUT;
  wire fifo16_READ_OUTPUT;
  wire fifo17_READ_OUTPUT;
  wire fifo18_READ_OUTPUT;
  wire fifo19_READ_OUTPUT;
  wire fifo20_READ_OUTPUT;
  wire fifo21_READ_OUTPUT;
  wire fifo22_READ_OUTPUT;
  wire fifo23_READ_OUTPUT;
  wire fifo24_READ_OUTPUT;
  wire [7:0] writeAddr_GET_OUTPUT;
  wire unnamedunary34984USEDMULTIPLEunary;assign unnamedunary34984USEDMULTIPLEunary = {(~{(writeAddr_GET_OUTPUT==readAddr_GET_OUTPUT)})}; 
  always @(posedge CLK) begin if(unnamedunary34984USEDMULTIPLEunary == 1'b0 && popFront_valid==1'b1 && CE_pop==1'b1) begin $display("%s: attempting to pop from an empty fifo",INSTANCE_NAME);$finish();  end end
  wire [7:0] readAddr_SETBY_OUTPUT;
  assign popFront = {fifo24_READ_OUTPUT,fifo23_READ_OUTPUT,fifo22_READ_OUTPUT,fifo21_READ_OUTPUT,fifo20_READ_OUTPUT,fifo19_READ_OUTPUT,fifo18_READ_OUTPUT,fifo17_READ_OUTPUT,fifo16_READ_OUTPUT,fifo15_READ_OUTPUT,fifo14_READ_OUTPUT,fifo13_READ_OUTPUT,fifo12_READ_OUTPUT,fifo11_READ_OUTPUT,fifo10_READ_OUTPUT,fifo9_READ_OUTPUT,fifo8_READ_OUTPUT,fifo7_READ_OUTPUT,fifo6_READ_OUTPUT,fifo5_READ_OUTPUT,fifo4_READ_OUTPUT,fifo3_READ_OUTPUT,fifo2_READ_OUTPUT,fifo1_READ_OUTPUT};
  wire [7:0] unnamedselect34975USEDMULTIPLEselect;assign unnamedselect34975USEDMULTIPLEselect = (({((writeAddr_GET_OUTPUT)<(readAddr_GET_OUTPUT))})?({({((8'd128)-readAddr_GET_OUTPUT)}+writeAddr_GET_OUTPUT)}):({(writeAddr_GET_OUTPUT-readAddr_GET_OUTPUT)})); 
  assign size = unnamedselect34975USEDMULTIPLEselect;
  reg readyReg;
    always @ (posedge CLK) begin readyReg <= {((unnamedselect34975USEDMULTIPLEselect)<((8'd125)))}; end
  assign ready = readyReg;
  always @(posedge CLK) begin if({((unnamedselect34975USEDMULTIPLEselect)<((8'd126)))} == 1'b0 && pushBack_valid==1'b1 && CE_push==1'b1) begin $display("%s: attempting to push to a full fifo",INSTANCE_NAME);$finish();  end end
  wire [7:0] writeAddr_SETBY_OUTPUT;
  wire [6:0] unnamedcast34992USEDMULTIPLEcast;assign unnamedcast34992USEDMULTIPLEcast = writeAddr_GET_OUTPUT[6:0]; 
  assign hasData = unnamedunary34984USEDMULTIPLEunary;
  // function: popFront pure=false delay=0
  // function: size pure=true delay=0
  // function: pushBackReset pure=false delay=0
  // function: ready pure=true delay=0
  // function: pushBack pure=false delay=0
  // function: popFrontReset pure=false delay=0
  // function: hasData pure=true delay=0
  RegBy_incif_wrapuint8_127_incnil_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_writeAddr"})) writeAddr(.CLK(CLK), .set_valid(pushBackReset_valid), .CE(CE_push), .set_inp((8'd0)), .setby_valid(pushBack_valid), .setby_inp((1'd1)), .SETBY_OUTPUT(writeAddr_SETBY_OUTPUT), .GET_OUTPUT(writeAddr_GET_OUTPUT));
  RegBy_incif_wrapuint8_127_incnil_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_readAddr"})) readAddr(.CLK(CLK), .set_valid(popFrontReset_valid), .CE(CE_pop), .set_inp((8'd0)), .setby_valid(popFront_valid), .setby_inp((1'd1)), .SETBY_OUTPUT(readAddr_SETBY_OUTPUT), .GET_OUTPUT(readAddr_GET_OUTPUT));
  wire [7:0] fifo1_writeInput = {pushBack_input[0:0],unnamedcast34992USEDMULTIPLEcast};
wire fifo1_writeOut;
RAM128X1D fifo1  (
  .WCLK(CLK),
  .D(fifo1_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo1_writeOut),
  .DPO(fifo1_READ_OUTPUT),
  .A(fifo1_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo2_writeInput = {pushBack_input[1:1],unnamedcast34992USEDMULTIPLEcast};
wire fifo2_writeOut;
RAM128X1D fifo2  (
  .WCLK(CLK),
  .D(fifo2_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo2_writeOut),
  .DPO(fifo2_READ_OUTPUT),
  .A(fifo2_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo3_writeInput = {pushBack_input[2:2],unnamedcast34992USEDMULTIPLEcast};
wire fifo3_writeOut;
RAM128X1D fifo3  (
  .WCLK(CLK),
  .D(fifo3_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo3_writeOut),
  .DPO(fifo3_READ_OUTPUT),
  .A(fifo3_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo4_writeInput = {pushBack_input[3:3],unnamedcast34992USEDMULTIPLEcast};
wire fifo4_writeOut;
RAM128X1D fifo4  (
  .WCLK(CLK),
  .D(fifo4_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo4_writeOut),
  .DPO(fifo4_READ_OUTPUT),
  .A(fifo4_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo5_writeInput = {pushBack_input[4:4],unnamedcast34992USEDMULTIPLEcast};
wire fifo5_writeOut;
RAM128X1D fifo5  (
  .WCLK(CLK),
  .D(fifo5_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo5_writeOut),
  .DPO(fifo5_READ_OUTPUT),
  .A(fifo5_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo6_writeInput = {pushBack_input[5:5],unnamedcast34992USEDMULTIPLEcast};
wire fifo6_writeOut;
RAM128X1D fifo6  (
  .WCLK(CLK),
  .D(fifo6_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo6_writeOut),
  .DPO(fifo6_READ_OUTPUT),
  .A(fifo6_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo7_writeInput = {pushBack_input[6:6],unnamedcast34992USEDMULTIPLEcast};
wire fifo7_writeOut;
RAM128X1D fifo7  (
  .WCLK(CLK),
  .D(fifo7_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo7_writeOut),
  .DPO(fifo7_READ_OUTPUT),
  .A(fifo7_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo8_writeInput = {pushBack_input[7:7],unnamedcast34992USEDMULTIPLEcast};
wire fifo8_writeOut;
RAM128X1D fifo8  (
  .WCLK(CLK),
  .D(fifo8_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo8_writeOut),
  .DPO(fifo8_READ_OUTPUT),
  .A(fifo8_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo9_writeInput = {pushBack_input[8:8],unnamedcast34992USEDMULTIPLEcast};
wire fifo9_writeOut;
RAM128X1D fifo9  (
  .WCLK(CLK),
  .D(fifo9_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo9_writeOut),
  .DPO(fifo9_READ_OUTPUT),
  .A(fifo9_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo10_writeInput = {pushBack_input[9:9],unnamedcast34992USEDMULTIPLEcast};
wire fifo10_writeOut;
RAM128X1D fifo10  (
  .WCLK(CLK),
  .D(fifo10_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo10_writeOut),
  .DPO(fifo10_READ_OUTPUT),
  .A(fifo10_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo11_writeInput = {pushBack_input[10:10],unnamedcast34992USEDMULTIPLEcast};
wire fifo11_writeOut;
RAM128X1D fifo11  (
  .WCLK(CLK),
  .D(fifo11_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo11_writeOut),
  .DPO(fifo11_READ_OUTPUT),
  .A(fifo11_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo12_writeInput = {pushBack_input[11:11],unnamedcast34992USEDMULTIPLEcast};
wire fifo12_writeOut;
RAM128X1D fifo12  (
  .WCLK(CLK),
  .D(fifo12_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo12_writeOut),
  .DPO(fifo12_READ_OUTPUT),
  .A(fifo12_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo13_writeInput = {pushBack_input[12:12],unnamedcast34992USEDMULTIPLEcast};
wire fifo13_writeOut;
RAM128X1D fifo13  (
  .WCLK(CLK),
  .D(fifo13_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo13_writeOut),
  .DPO(fifo13_READ_OUTPUT),
  .A(fifo13_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo14_writeInput = {pushBack_input[13:13],unnamedcast34992USEDMULTIPLEcast};
wire fifo14_writeOut;
RAM128X1D fifo14  (
  .WCLK(CLK),
  .D(fifo14_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo14_writeOut),
  .DPO(fifo14_READ_OUTPUT),
  .A(fifo14_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo15_writeInput = {pushBack_input[14:14],unnamedcast34992USEDMULTIPLEcast};
wire fifo15_writeOut;
RAM128X1D fifo15  (
  .WCLK(CLK),
  .D(fifo15_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo15_writeOut),
  .DPO(fifo15_READ_OUTPUT),
  .A(fifo15_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo16_writeInput = {pushBack_input[15:15],unnamedcast34992USEDMULTIPLEcast};
wire fifo16_writeOut;
RAM128X1D fifo16  (
  .WCLK(CLK),
  .D(fifo16_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo16_writeOut),
  .DPO(fifo16_READ_OUTPUT),
  .A(fifo16_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo17_writeInput = {pushBack_input[16:16],unnamedcast34992USEDMULTIPLEcast};
wire fifo17_writeOut;
RAM128X1D fifo17  (
  .WCLK(CLK),
  .D(fifo17_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo17_writeOut),
  .DPO(fifo17_READ_OUTPUT),
  .A(fifo17_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo18_writeInput = {pushBack_input[17:17],unnamedcast34992USEDMULTIPLEcast};
wire fifo18_writeOut;
RAM128X1D fifo18  (
  .WCLK(CLK),
  .D(fifo18_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo18_writeOut),
  .DPO(fifo18_READ_OUTPUT),
  .A(fifo18_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo19_writeInput = {pushBack_input[18:18],unnamedcast34992USEDMULTIPLEcast};
wire fifo19_writeOut;
RAM128X1D fifo19  (
  .WCLK(CLK),
  .D(fifo19_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo19_writeOut),
  .DPO(fifo19_READ_OUTPUT),
  .A(fifo19_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo20_writeInput = {pushBack_input[19:19],unnamedcast34992USEDMULTIPLEcast};
wire fifo20_writeOut;
RAM128X1D fifo20  (
  .WCLK(CLK),
  .D(fifo20_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo20_writeOut),
  .DPO(fifo20_READ_OUTPUT),
  .A(fifo20_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo21_writeInput = {pushBack_input[20:20],unnamedcast34992USEDMULTIPLEcast};
wire fifo21_writeOut;
RAM128X1D fifo21  (
  .WCLK(CLK),
  .D(fifo21_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo21_writeOut),
  .DPO(fifo21_READ_OUTPUT),
  .A(fifo21_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo22_writeInput = {pushBack_input[21:21],unnamedcast34992USEDMULTIPLEcast};
wire fifo22_writeOut;
RAM128X1D fifo22  (
  .WCLK(CLK),
  .D(fifo22_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo22_writeOut),
  .DPO(fifo22_READ_OUTPUT),
  .A(fifo22_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo23_writeInput = {pushBack_input[22:22],unnamedcast34992USEDMULTIPLEcast};
wire fifo23_writeOut;
RAM128X1D fifo23  (
  .WCLK(CLK),
  .D(fifo23_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo23_writeOut),
  .DPO(fifo23_READ_OUTPUT),
  .A(fifo23_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

  wire [7:0] fifo24_writeInput = {pushBack_input[23:23],unnamedcast34992USEDMULTIPLEcast};
wire fifo24_writeOut;
RAM128X1D fifo24  (
  .WCLK(CLK),
  .D(fifo24_writeInput[7]),
  .WE(pushBack_valid && CE_push),
  .SPO(fifo24_writeOut),
  .DPO(fifo24_READ_OUTPUT),
  .A(fifo24_writeInput[6:0]),
  .DPRA(unnamedcast35117USEDMULTIPLEcast));

endmodule

module fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384(input CLK, input load_valid, input load_CE, output [24:0] load_output, input store_reset_valid, input store_CE, output store_ready, input load_reset_valid, input store_valid, input [23:0] store_input);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(load_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_reset_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(load_reset_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store'", INSTANCE_NAME);  end end
  wire FIFO_hasData;
  wire [23:0] FIFO_popFront;
  assign load_output = {FIFO_hasData,FIFO_popFront};
  wire FIFO_ready;
  assign store_ready = FIFO_ready;
  // function: load pure=false delay=0
  // function: store_reset pure=false delay=0
  // function: store_ready pure=true delay=0
  // function: load_reset pure=false delay=0
  // function: store pure=false delay=0
  fifo__uint8_uint16__128 #(.INSTANCE_NAME({INSTANCE_NAME,"_FIFO"})) FIFO(.CLK(CLK), .popFront_valid({(FIFO_hasData&&load_valid)}), .CE_pop(load_CE), .popFront(FIFO_popFront), .size(FIFO_size), .pushBackReset_valid(store_reset_valid), .CE_push(store_CE), .ready(FIFO_ready), .pushBack_valid(store_valid), .pushBack_input(store_input), .popFrontReset_valid(load_reset_valid), .hasData(FIFO_hasData));
endmodule

module LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384(input CLK, input load_valid, input load_CE, input load_input, output [24:0] load_output, input store_reset_valid, input store_CE, output store_ready, output load_ready, input load_reset, input store_valid, input [23:0] store_input);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(load_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_reset_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(load_reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store'", INSTANCE_NAME);  end end
  wire unnamedcast35616USEDMULTIPLEcast;assign unnamedcast35616USEDMULTIPLEcast = load_input; 
  wire [24:0] LiftDecimate_load_output;
  reg [23:0] unnamedcast35619_delay1_validunnamednull0_CEload_CE;  always @ (posedge CLK) begin if (load_CE) begin unnamedcast35619_delay1_validunnamednull0_CEload_CE <= (LiftDecimate_load_output[23:0]); end end
  reg unnamedbinop35624_delay1_validunnamednull0_CEload_CE;  always @ (posedge CLK) begin if (load_CE) begin unnamedbinop35624_delay1_validunnamednull0_CEload_CE <= {((LiftDecimate_load_output[24])&&unnamedcast35616USEDMULTIPLEcast)}; end end
  assign load_output = {unnamedbinop35624_delay1_validunnamednull0_CEload_CE,unnamedcast35619_delay1_validunnamednull0_CEload_CE};
  wire LiftDecimate_store_ready;
  assign store_ready = LiftDecimate_store_ready;
  assign load_ready = (1'd1);
  // function: load pure=false delay=1
  // function: store_reset pure=false delay=0
  // function: store_ready pure=true delay=0
  // function: load_ready pure=true delay=0
  // function: load_reset pure=false delay=0
  // function: store pure=false delay=0
  fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384 #(.INSTANCE_NAME({INSTANCE_NAME,"_LiftDecimate"})) LiftDecimate(.CLK(CLK), .load_valid({(unnamedcast35616USEDMULTIPLEcast&&load_valid)}), .load_CE(load_CE), .load_output(LiftDecimate_load_output), .store_reset_valid(store_reset_valid), .store_CE(store_CE), .store_ready(LiftDecimate_store_ready), .load_reset_valid(load_reset), .store_valid(store_valid), .store_input(store_input));
endmodule

module RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384(input CLK, input load_valid, input load_CE, input load_input, output [24:0] load_output, input store_reset, input CE, output store_ready, output load_ready, input load_reset, input store_valid, input [24:0] store_input, output store_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(load_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(load_reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'load_reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(store_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'store'", INSTANCE_NAME);  end end
  wire [24:0] RunIffReady_load_output;
  assign load_output = RunIffReady_load_output;
  wire RunIffReady_store_ready;
  assign store_ready = RunIffReady_store_ready;
  wire RunIffReady_load_ready;
  assign load_ready = RunIffReady_load_ready;
  wire unnamedbinop35695USEDMULTIPLEbinop;assign unnamedbinop35695USEDMULTIPLEbinop = {({(RunIffReady_store_ready&&(store_input[24]))}&&store_valid)}; 
  assign store_output = {unnamedbinop35695USEDMULTIPLEbinop};
  // function: load pure=false delay=1
  // function: store_reset pure=false delay=0
  // function: store_ready pure=true delay=0
  // function: load_ready pure=true delay=0
  // function: load_reset pure=false delay=0
  // function: store pure=false delay=0
  LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384 #(.INSTANCE_NAME({INSTANCE_NAME,"_RunIffReady"})) RunIffReady(.CLK(CLK), .load_valid(load_valid), .load_CE(load_CE), .load_input(load_input), .load_output(RunIffReady_load_output), .store_reset_valid(store_reset), .store_CE(CE), .store_ready(RunIffReady_store_ready), .load_ready(RunIffReady_load_ready), .load_reset(load_reset), .store_valid(unnamedbinop35695USEDMULTIPLEbinop), .store_input((store_input[23:0])));
endmodule

module LiftHandshake_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384(input CLK, input load_input, output [24:0] load_output, input store_reset, input store_ready_downstream, output store_ready, input load_ready_downstream, output load_ready, input load_reset, input [24:0] store_input, output store_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire unnamedunary35732USEDMULTIPLEunary;assign unnamedunary35732USEDMULTIPLEunary = {(~load_reset)}; 
  wire unnamedbinop35731USEDMULTIPLEbinop;assign unnamedbinop35731USEDMULTIPLEbinop = {(load_reset||load_ready_downstream)}; 
  wire [24:0] inner_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384_load_output;
  wire load_validBitDelay_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384_pushPop_out;
  wire [24:0] unnamedtuple35742USEDMULTIPLEtuple;assign unnamedtuple35742USEDMULTIPLEtuple = {{((inner_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384_load_output[24])&&load_validBitDelay_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384_pushPop_out)},(inner_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384_load_output[23:0])}; 
  always @(posedge CLK) begin if({(~{((unnamedtuple35742USEDMULTIPLEtuple[24])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: output valid bit should not be X!",INSTANCE_NAME); end end
  always @(posedge CLK) begin if({(~{(load_input===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign load_output = unnamedtuple35742USEDMULTIPLEtuple;
  wire unnamedbinop35760USEDMULTIPLEbinop;assign unnamedbinop35760USEDMULTIPLEbinop = {(store_reset||store_ready_downstream)}; 
  wire inner_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384_store_ready;
  assign store_ready = {(inner_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384_store_ready&&store_ready_downstream)};
  wire inner_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384_load_ready;
  assign load_ready = {(inner_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384_load_ready&&load_ready_downstream)};
  wire unnamedunary35761USEDMULTIPLEunary;assign unnamedunary35761USEDMULTIPLEunary = {(~store_reset)}; 
  wire [0:0] inner_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384_store_output;
  wire store_validBitDelay_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384_pushPop_out;
  wire [0:0] unnamedtuple35771USEDMULTIPLEtuple;assign unnamedtuple35771USEDMULTIPLEtuple = {{(inner_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384_store_output&&store_validBitDelay_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384_pushPop_out)}}; 
  always @(posedge CLK) begin if({(~{(unnamedtuple35771USEDMULTIPLEtuple===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: output valid bit should not be X!",INSTANCE_NAME); end end
  always @(posedge CLK) begin if({(~{((store_input[24])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign store_output = unnamedtuple35771USEDMULTIPLEtuple;
  // function: load pure=false ONLY WIRE
  // function: store_reset pure=false ONLY WIRE
  // function: store_ready pure=true ONLY WIRE
  // function: load_ready pure=true ONLY WIRE
  // function: load_reset pure=false ONLY WIRE
  // function: store pure=false ONLY WIRE
  RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384 #(.INSTANCE_NAME({INSTANCE_NAME,"_inner_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384"})) inner_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384(.CLK(CLK), .load_valid(unnamedunary35732USEDMULTIPLEunary), .load_CE(unnamedbinop35731USEDMULTIPLEbinop), .load_input(load_input), .load_output(inner_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384_load_output), .store_reset(store_reset), .CE(unnamedbinop35760USEDMULTIPLEbinop), .store_ready(inner_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384_store_ready), .load_ready(inner_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384_load_ready), .load_reset(load_reset), .store_valid(unnamedunary35761USEDMULTIPLEunary), .store_input(store_input), .store_output(inner_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384_store_output));
  ShiftRegister_1_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_load_validBitDelay_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384"})) load_validBitDelay_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384(.CLK(CLK), .pushPop_valid(unnamedunary35732USEDMULTIPLEunary), .CE(unnamedbinop35731USEDMULTIPLEbinop), .sr_input((1'd1)), .pushPop_out(load_validBitDelay_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384_pushPop_out), .reset(load_reset));
  ShiftRegister_0_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_store_validBitDelay_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384"})) store_validBitDelay_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384(.CLK(CLK), .CE(unnamedbinop35760USEDMULTIPLEbinop), .sr_input((1'd1)), .pushPop_out(store_validBitDelay_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384_pushPop_out));
endmodule

module ShiftRegister_4_CEtrue_TY1(input CLK, input pushPop_valid, input CE, input sr_input, output pushPop_out, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'pushPop'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  reg SR4;
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR1' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR1' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR1' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate35935USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate35935USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(sr_input):((1'd0)))}; 
  reg SR1;  always @ (posedge CLK) begin if ((unnamedcallArbitrate35935USEDMULTIPLEcallArbitrate[1]) && CE) begin SR1 <= (unnamedcallArbitrate35935USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR2' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR2' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR2' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate35941USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate35941USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR1):((1'd0)))}; 
  reg SR2;  always @ (posedge CLK) begin if ((unnamedcallArbitrate35941USEDMULTIPLEcallArbitrate[1]) && CE) begin SR2 <= (unnamedcallArbitrate35941USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR3' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR3' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR3' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate35947USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate35947USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR2):((1'd0)))}; 
  reg SR3;  always @ (posedge CLK) begin if ((unnamedcallArbitrate35947USEDMULTIPLEcallArbitrate[1]) && CE) begin SR3 <= (unnamedcallArbitrate35947USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR4' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR4' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR4' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate35953USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate35953USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR3):((1'd0)))}; 
    always @ (posedge CLK) begin if ((unnamedcallArbitrate35953USEDMULTIPLEcallArbitrate[1]) && CE) begin SR4 <= (unnamedcallArbitrate35953USEDMULTIPLEcallArbitrate[0]); end end
  assign pushPop_out = SR4;
  // function: pushPop pure=false delay=0
  // function: reset pure=false delay=0
endmodule

module displayOutput(input CLK, input process_CE, input [23:0] inp, output [31:0] process_output);
parameter INSTANCE_NAME="INST";
  reg unnamedbinop35825_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop35825_delay1_validunnamednull0_CEprocess_CE <= {(((inp[23:8]))<((16'd2144)))}; end end
  reg unnamedbinop35825_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop35825_delay2_validunnamednull0_CEprocess_CE <= unnamedbinop35825_delay1_validunnamednull0_CEprocess_CE; end end
  reg unnamedbinop35825_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop35825_delay3_validunnamednull0_CEprocess_CE <= unnamedbinop35825_delay2_validunnamednull0_CEprocess_CE; end end
  reg [31:0] unnamedcast35820_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast35820_delay1_validunnamednull0_CEprocess_CE <= {{(8'd0),(8'd0),(8'd0),(8'd0)}}; end end
  reg [31:0] unnamedcast35820_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast35820_delay2_validunnamednull0_CEprocess_CE <= unnamedcast35820_delay1_validunnamednull0_CEprocess_CE; end end
  reg [31:0] unnamedcast35820_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast35820_delay3_validunnamednull0_CEprocess_CE <= unnamedcast35820_delay2_validunnamednull0_CEprocess_CE; end end
  reg [7:0] unnamedbinop35797_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop35797_delay1_validunnamednull0_CEprocess_CE <= {((inp[7:0])-(8'd60))}; end end
  reg [7:0] unnamedcast35799_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast35799_delay1_validunnamednull0_CEprocess_CE <= (8'd4); end end
  reg [7:0] unnamedbinop35800_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop35800_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop35797_delay1_validunnamednull0_CEprocess_CE<<<unnamedcast35799_delay1_validunnamednull0_CEprocess_CE)}; end end
  reg [7:0] unnamedbinop35800_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop35800_delay2_validunnamednull0_CEprocess_CE <= unnamedbinop35800_delay1_validunnamednull0_CEprocess_CE; end end
  reg [7:0] unnamedcast35808_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast35808_delay1_validunnamednull0_CEprocess_CE <= (8'd16); end end
  reg [7:0] unnamedbinop35809_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop35809_delay1_validunnamednull0_CEprocess_CE <= {(unnamedcast35808_delay1_validunnamednull0_CEprocess_CE-unnamedbinop35797_delay1_validunnamednull0_CEprocess_CE)}; end end
  reg [7:0] unnamedcast35799_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast35799_delay2_validunnamednull0_CEprocess_CE <= unnamedcast35799_delay1_validunnamednull0_CEprocess_CE; end end
  reg [7:0] unnamedbinop35812_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop35812_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop35809_delay1_validunnamednull0_CEprocess_CE<<<unnamedcast35799_delay2_validunnamednull0_CEprocess_CE)}; end end
  reg [31:0] unnamedselect35826_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedselect35826_delay1_validunnamednull0_CEprocess_CE <= ((unnamedbinop35825_delay3_validunnamednull0_CEprocess_CE)?(unnamedcast35820_delay3_validunnamednull0_CEprocess_CE):({{(8'd0),unnamedbinop35812_delay1_validunnamednull0_CEprocess_CE,(8'd128),unnamedbinop35800_delay2_validunnamednull0_CEprocess_CE}})); end end
  assign process_output = unnamedselect35826_delay1_validunnamednull0_CEprocess_CE;
  // function: process pure=true delay=4
endmodule

module MakeHandshake_displayOutput(input CLK, input ready_downstream, output ready, input reset, input [24:0] process_input, output [32:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  assign ready = ready_downstream;
  wire unnamedbinop35965USEDMULTIPLEbinop;assign unnamedbinop35965USEDMULTIPLEbinop = {(ready_downstream||reset)}; 
  wire unnamedcast35973USEDMULTIPLEcast;assign unnamedcast35973USEDMULTIPLEcast = (process_input[24]); 
  wire [31:0] inner_process_output;
  wire validBitDelay_displayOutput_pushPop_out;
  always @(posedge CLK) begin if({(~{(unnamedcast35973USEDMULTIPLEcast===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: MakeHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = {validBitDelay_displayOutput_pushPop_out,inner_process_output};
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  ShiftRegister_4_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_validBitDelay_displayOutput"})) validBitDelay_displayOutput(.CLK(CLK), .pushPop_valid({(~reset)}), .CE(unnamedbinop35965USEDMULTIPLEbinop), .sr_input(unnamedcast35973USEDMULTIPLEcast), .pushPop_out(validBitDelay_displayOutput_pushPop_out), .reset(reset));
  displayOutput #(.INSTANCE_NAME({INSTANCE_NAME,"_inner"})) inner(.CLK(CLK), .process_CE(unnamedbinop35965USEDMULTIPLEbinop), .inp((process_input[23:0])), .process_output(inner_process_output));
endmodule

module incif_wrapuint16_830_inc1(input CLK, input CE, input [16:0] process_input, output [15:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] unnamedcast308USEDMULTIPLEcast;assign unnamedcast308USEDMULTIPLEcast = (process_input[15:0]); 
  assign process_output = (((process_input[16]))?((({(unnamedcast308USEDMULTIPLEcast==(16'd830))})?((16'd0)):({(unnamedcast308USEDMULTIPLEcast+(16'd1))}))):(unnamedcast308USEDMULTIPLEcast));
  // function: process pure=true delay=0
endmodule

module RegBy_incif_wrapuint16_830_inc1_CEtrue_init0(input CLK, input set_valid, input CE, input [15:0] set_inp, input setby_valid, input setby_inp, output [15:0] SETBY_OUTPUT, output [15:0] GET_OUTPUT);
parameter INSTANCE_NAME="INST";
  reg [15:0] R = 16'd0;
  wire [15:0] regby_inner_process_output;
  always @(posedge CLK) begin if(set_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(setby_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,set_valid})+({4'b0,setby_valid})) > 5'd1) begin $display("error, function 'set' on instance 'R' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [16:0] unnamedcallArbitrate359USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate359USEDMULTIPLEcallArbitrate = {(set_valid||setby_valid),((set_valid)?(set_inp):(regby_inner_process_output))}; 
    always @ (posedge CLK) begin if ((unnamedcallArbitrate359USEDMULTIPLEcallArbitrate[16]) && CE) begin R <= (unnamedcallArbitrate359USEDMULTIPLEcallArbitrate[15:0]); end end
  assign SETBY_OUTPUT = regby_inner_process_output;
  assign GET_OUTPUT = R;
  // function: set pure=false ONLY WIRE
  // function: setby pure=false ONLY WIRE
  // function: get pure=true ONLY WIRE
  incif_wrapuint16_830_inc1 #(.INSTANCE_NAME({INSTANCE_NAME,"_regby_inner"})) regby_inner(.CLK(CLK), .CE(CE), .process_input({setby_inp,R}), .process_output(regby_inner_process_output));
endmodule

module incif_wrapuint16_494_incnil(input CLK, input CE, input [16:0] process_input, output [15:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] unnamedcast366USEDMULTIPLEcast;assign unnamedcast366USEDMULTIPLEcast = (process_input[15:0]); 
  assign process_output = (((process_input[16]))?((({(unnamedcast366USEDMULTIPLEcast==(16'd494))})?((16'd0)):({(unnamedcast366USEDMULTIPLEcast+(16'd1))}))):(unnamedcast366USEDMULTIPLEcast));
  // function: process pure=true delay=0
endmodule

module RegBy_incif_wrapuint16_494_incnil_CEtrue_init0(input CLK, input set_valid, input CE, input [15:0] set_inp, input setby_valid, input setby_inp, output [15:0] SETBY_OUTPUT, output [15:0] GET_OUTPUT);
parameter INSTANCE_NAME="INST";
  reg [15:0] R = 16'd0;
  wire [15:0] regby_inner_process_output;
  always @(posedge CLK) begin if(set_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(setby_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,set_valid})+({4'b0,setby_valid})) > 5'd1) begin $display("error, function 'set' on instance 'R' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [16:0] unnamedcallArbitrate417USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate417USEDMULTIPLEcallArbitrate = {(set_valid||setby_valid),((set_valid)?(set_inp):(regby_inner_process_output))}; 
    always @ (posedge CLK) begin if ((unnamedcallArbitrate417USEDMULTIPLEcallArbitrate[16]) && CE) begin R <= (unnamedcallArbitrate417USEDMULTIPLEcallArbitrate[15:0]); end end
  assign SETBY_OUTPUT = regby_inner_process_output;
  assign GET_OUTPUT = R;
  // function: set pure=false ONLY WIRE
  // function: setby pure=false ONLY WIRE
  // function: get pure=true ONLY WIRE
  incif_wrapuint16_494_incnil #(.INSTANCE_NAME({INSTANCE_NAME,"_regby_inner"})) regby_inner(.CLK(CLK), .CE(CE), .process_input({setby_inp,R}), .process_output(regby_inner_process_output));
endmodule

module PosSeq_W831_H495_T1(input CLK, input process_valid, input CE, output [31:0] process_output, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  wire [15:0] posX_posSeq_GET_OUTPUT;
  wire [15:0] posY_posSeq_GET_OUTPUT;
  wire [15:0] posX_posSeq_SETBY_OUTPUT;
  wire [15:0] posY_posSeq_SETBY_OUTPUT;
  assign process_output = {{posY_posSeq_GET_OUTPUT,posX_posSeq_GET_OUTPUT}};
  // function: process pure=false delay=0
  // function: reset pure=false delay=0
  RegBy_incif_wrapuint16_830_inc1_CEtrue_init0 #(.INSTANCE_NAME({INSTANCE_NAME,"_posX_posSeq"})) posX_posSeq(.CLK(CLK), .set_valid(reset), .CE(CE), .set_inp((16'd0)), .setby_valid(process_valid), .setby_inp((1'd1)), .SETBY_OUTPUT(posX_posSeq_SETBY_OUTPUT), .GET_OUTPUT(posX_posSeq_GET_OUTPUT));
  RegBy_incif_wrapuint16_494_incnil_CEtrue_init0 #(.INSTANCE_NAME({INSTANCE_NAME,"_posY_posSeq"})) posY_posSeq(.CLK(CLK), .set_valid(reset), .CE(CE), .set_inp((16'd0)), .setby_valid(process_valid), .setby_inp({(posX_posSeq_GET_OUTPUT==(16'd830))}), .SETBY_OUTPUT(posY_posSeq_SETBY_OUTPUT), .GET_OUTPUT(posY_posSeq_GET_OUTPUT));
endmodule

module CropSeq_uint8_4_1__W831_H495_T1(input CLK, input process_CE, input [63:0] process_input, output [32:0] process_output);
parameter INSTANCE_NAME="INST";
  reg [31:0] unnamedcast35978_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast35978_delay1_validunnamednull0_CEprocess_CE <= (process_input[63:32]); end end
  reg [31:0] unnamedcast35978_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast35978_delay2_validunnamednull0_CEprocess_CE <= unnamedcast35978_delay1_validunnamednull0_CEprocess_CE; end end
  reg [31:0] unnamedcast35978_delay3_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast35978_delay3_validunnamednull0_CEprocess_CE <= unnamedcast35978_delay2_validunnamednull0_CEprocess_CE; end end
  wire [31:0] unnamedcast35980;assign unnamedcast35980 = (process_input[31:0]);  // wire for array index
  wire [31:0] unnamedcast35982USEDMULTIPLEcast;assign unnamedcast35982USEDMULTIPLEcast = ({unnamedcast35980[31:0]}); 
  wire [15:0] unnamedcast35984USEDMULTIPLEcast;assign unnamedcast35984USEDMULTIPLEcast = (unnamedcast35982USEDMULTIPLEcast[15:0]); 
  reg unnamedbinop35996_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop35996_delay1_validunnamednull0_CEprocess_CE <= {((unnamedcast35984USEDMULTIPLEcast)>=((16'd191)))}; end end
  wire [15:0] unnamedcast35990USEDMULTIPLEcast;assign unnamedcast35990USEDMULTIPLEcast = (unnamedcast35982USEDMULTIPLEcast[31:16]); 
  reg unnamedbinop35998_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop35998_delay1_validunnamednull0_CEprocess_CE <= {((unnamedcast35990USEDMULTIPLEcast)>=((16'd15)))}; end end
  reg unnamedbinop35999_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop35999_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop35996_delay1_validunnamednull0_CEprocess_CE&&unnamedbinop35998_delay1_validunnamednull0_CEprocess_CE)}; end end
  reg unnamedbinop36001_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop36001_delay1_validunnamednull0_CEprocess_CE <= {((unnamedcast35984USEDMULTIPLEcast)<((16'd831)))}; end end
  reg unnamedbinop36003_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop36003_delay1_validunnamednull0_CEprocess_CE <= {((unnamedcast35990USEDMULTIPLEcast)<((16'd495)))}; end end
  reg unnamedbinop36004_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop36004_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop36001_delay1_validunnamednull0_CEprocess_CE&&unnamedbinop36003_delay1_validunnamednull0_CEprocess_CE)}; end end
  reg unnamedbinop36005_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop36005_delay1_validunnamednull0_CEprocess_CE <= {(unnamedbinop35999_delay1_validunnamednull0_CEprocess_CE&&unnamedbinop36004_delay1_validunnamednull0_CEprocess_CE)}; end end
  assign process_output = {unnamedbinop36005_delay1_validunnamednull0_CEprocess_CE,unnamedcast35978_delay3_validunnamednull0_CEprocess_CE};
  // function: process pure=true delay=3
endmodule

module liftXYSeq_lift_CropSeq_uint8_4_1__W831_H495_T1(input CLK, input process_valid, input CE, input [31:0] process_input, output [32:0] process_output, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  wire [31:0] p_process_output;
  wire [32:0] m_process_output;
  assign process_output = m_process_output;
  // function: process pure=false delay=3
  // function: reset pure=false delay=0
  PosSeq_W831_H495_T1 #(.INSTANCE_NAME({INSTANCE_NAME,"_p"})) p(.CLK(CLK), .process_valid(process_valid), .CE(CE), .process_output(p_process_output), .reset(reset));
  CropSeq_uint8_4_1__W831_H495_T1 #(.INSTANCE_NAME({INSTANCE_NAME,"_m"})) m(.CLK(CLK), .process_CE(CE), .process_input({process_input,p_process_output}), .process_output(m_process_output));
endmodule

module LiftDecimate_liftXYSeq_lift_CropSeq_uint8_4_1__W831_H495_T1(input CLK, output ready, input reset, input CE, input process_valid, input [32:0] process_input, output [32:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  assign ready = (1'd1);
  wire unnamedcast36120USEDMULTIPLEcast;assign unnamedcast36120USEDMULTIPLEcast = (process_input[32]); 
  wire [32:0] LiftDecimate_process_output;
  reg [31:0] unnamedcast36123_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast36123_delay1_validunnamednull0_CECE <= (LiftDecimate_process_output[31:0]); end end
  reg unnamedcast36120_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast36120_delay1_validunnamednull0_CECE <= unnamedcast36120USEDMULTIPLEcast; end end
  reg unnamedcast36120_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast36120_delay2_validunnamednull0_CECE <= unnamedcast36120_delay1_validunnamednull0_CECE; end end
  reg unnamedcast36120_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast36120_delay3_validunnamednull0_CECE <= unnamedcast36120_delay2_validunnamednull0_CECE; end end
  reg unnamedbinop36128_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedbinop36128_delay1_validunnamednull0_CECE <= {((LiftDecimate_process_output[32])&&unnamedcast36120_delay3_validunnamednull0_CECE)}; end end
  assign process_output = {unnamedbinop36128_delay1_validunnamednull0_CECE,unnamedcast36123_delay1_validunnamednull0_CECE};
  // function: ready pure=true delay=0
  // function: reset pure=false delay=0
  // function: process pure=false delay=4
  liftXYSeq_lift_CropSeq_uint8_4_1__W831_H495_T1 #(.INSTANCE_NAME({INSTANCE_NAME,"_LiftDecimate"})) LiftDecimate(.CLK(CLK), .process_valid({(unnamedcast36120USEDMULTIPLEcast&&process_valid)}), .CE(CE), .process_input((process_input[31:0])), .process_output(LiftDecimate_process_output), .reset(reset));
endmodule

module LiftHandshake_LiftDecimate_liftXYSeq_lift_CropSeq_uint8_4_1__W831_H495_T1(input CLK, input ready_downstream, output ready, input reset, input [32:0] process_input, output [32:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire inner_LiftDecimate_liftXYSeq_lift_CropSeq_uint8_4_1__W831_H495_T1_ready;
  assign ready = {(inner_LiftDecimate_liftXYSeq_lift_CropSeq_uint8_4_1__W831_H495_T1_ready&&ready_downstream)};
  wire unnamedbinop36167USEDMULTIPLEbinop;assign unnamedbinop36167USEDMULTIPLEbinop = {(reset||ready_downstream)}; 
  wire unnamedunary36168USEDMULTIPLEunary;assign unnamedunary36168USEDMULTIPLEunary = {(~reset)}; 
  wire [32:0] inner_LiftDecimate_liftXYSeq_lift_CropSeq_uint8_4_1__W831_H495_T1_process_output;
  wire validBitDelay_LiftDecimate_liftXYSeq_lift_CropSeq_uint8_4_1__W831_H495_T1_pushPop_out;
  wire [32:0] unnamedtuple36178USEDMULTIPLEtuple;assign unnamedtuple36178USEDMULTIPLEtuple = {{((inner_LiftDecimate_liftXYSeq_lift_CropSeq_uint8_4_1__W831_H495_T1_process_output[32])&&validBitDelay_LiftDecimate_liftXYSeq_lift_CropSeq_uint8_4_1__W831_H495_T1_pushPop_out)},(inner_LiftDecimate_liftXYSeq_lift_CropSeq_uint8_4_1__W831_H495_T1_process_output[31:0])}; 
  always @(posedge CLK) begin if({(~{((unnamedtuple36178USEDMULTIPLEtuple[32])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: output valid bit should not be X!",INSTANCE_NAME); end end
  always @(posedge CLK) begin if({(~{((process_input[32])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = unnamedtuple36178USEDMULTIPLEtuple;
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  LiftDecimate_liftXYSeq_lift_CropSeq_uint8_4_1__W831_H495_T1 #(.INSTANCE_NAME({INSTANCE_NAME,"_inner_LiftDecimate_liftXYSeq_lift_CropSeq_uint8_4_1__W831_H495_T1"})) inner_LiftDecimate_liftXYSeq_lift_CropSeq_uint8_4_1__W831_H495_T1(.CLK(CLK), .ready(inner_LiftDecimate_liftXYSeq_lift_CropSeq_uint8_4_1__W831_H495_T1_ready), .reset(reset), .CE(unnamedbinop36167USEDMULTIPLEbinop), .process_valid(unnamedunary36168USEDMULTIPLEunary), .process_input(process_input), .process_output(inner_LiftDecimate_liftXYSeq_lift_CropSeq_uint8_4_1__W831_H495_T1_process_output));
  ShiftRegister_4_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_validBitDelay_LiftDecimate_liftXYSeq_lift_CropSeq_uint8_4_1__W831_H495_T1"})) validBitDelay_LiftDecimate_liftXYSeq_lift_CropSeq_uint8_4_1__W831_H495_T1(.CLK(CLK), .pushPop_valid(unnamedunary36168USEDMULTIPLEunary), .CE(unnamedbinop36167USEDMULTIPLEbinop), .sr_input((1'd1)), .pushPop_out(validBitDelay_LiftDecimate_liftXYSeq_lift_CropSeq_uint8_4_1__W831_H495_T1_pushPop_out), .reset(reset));
endmodule

module incif_wrapuint16_1_incnil(input CLK, input CE, input [16:0] process_input, output [15:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] unnamedcast36197USEDMULTIPLEcast;assign unnamedcast36197USEDMULTIPLEcast = (process_input[15:0]); 
  wire [15:0] unnamedcast36199USEDMULTIPLEcast;assign unnamedcast36199USEDMULTIPLEcast = (16'd1); 
  assign process_output = (((process_input[16]))?((({(unnamedcast36197USEDMULTIPLEcast==unnamedcast36199USEDMULTIPLEcast)})?((16'd0)):({(unnamedcast36197USEDMULTIPLEcast+unnamedcast36199USEDMULTIPLEcast)}))):(unnamedcast36197USEDMULTIPLEcast));
  // function: process pure=true delay=0
endmodule

module RegBy_incif_wrapuint16_1_incnil_CEtrue_initnil(input CLK, input set_valid, input CE, input [15:0] set_inp, input setby_valid, input setby_inp, output [15:0] SETBY_OUTPUT, output [15:0] GET_OUTPUT);
parameter INSTANCE_NAME="INST";
  reg [15:0] R;
  wire [15:0] regby_inner_process_output;
  always @(posedge CLK) begin if(set_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(setby_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,set_valid})+({4'b0,setby_valid})) > 5'd1) begin $display("error, function 'set' on instance 'R' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [16:0] unnamedcallArbitrate36248USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate36248USEDMULTIPLEcallArbitrate = {(set_valid||setby_valid),((set_valid)?(set_inp):(regby_inner_process_output))}; 
    always @ (posedge CLK) begin if ((unnamedcallArbitrate36248USEDMULTIPLEcallArbitrate[16]) && CE) begin R <= (unnamedcallArbitrate36248USEDMULTIPLEcallArbitrate[15:0]); end end
  assign SETBY_OUTPUT = regby_inner_process_output;
  assign GET_OUTPUT = R;
  // function: set pure=false ONLY WIRE
  // function: setby pure=false ONLY WIRE
  // function: get pure=true ONLY WIRE
  incif_wrapuint16_1_incnil #(.INSTANCE_NAME({INSTANCE_NAME,"_regby_inner"})) regby_inner(.CLK(CLK), .CE(CE), .process_input({setby_inp,R}), .process_output(regby_inner_process_output));
endmodule

module ChangeRate_uint8_4_1__from1_to2_H1(input CLK, output ready, input reset, input CE, input process_valid, input [31:0] process_input, output [64:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  assign ready = (1'd1);
  reg [31:0] process_input_delay1_validprocess_valid_CECE;  always @ (posedge CLK) begin if (process_valid && CE) begin process_input_delay1_validprocess_valid_CECE <= process_input; end end
  wire [15:0] phase_changerateup_GET_OUTPUT;
  wire [15:0] phase_changerateup_SETBY_OUTPUT;
  assign process_output = {{(phase_changerateup_GET_OUTPUT==(16'd1))},{({process_input[31:0]}),({process_input_delay1_validprocess_valid_CECE[31:0]})}};
  // function: ready pure=true delay=0
  // function: reset pure=false delay=0
  // function: process pure=false delay=0
  RegBy_incif_wrapuint16_1_incnil_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_phase_changerateup"})) phase_changerateup(.CLK(CLK), .set_valid(reset), .CE(CE), .set_inp((16'd0)), .setby_valid(process_valid), .setby_inp((1'd1)), .SETBY_OUTPUT(phase_changerateup_SETBY_OUTPUT), .GET_OUTPUT(phase_changerateup_GET_OUTPUT));
endmodule

module WaitOnInput_ChangeRate_uint8_4_1__from1_to2_H1(input CLK, output ready, input reset, input CE, input process_valid, input [32:0] process_input, output [64:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  wire WaitOnInput_inner_ready;
  assign ready = WaitOnInput_inner_ready;
  wire unnamedbinop36316USEDMULTIPLEbinop;assign unnamedbinop36316USEDMULTIPLEbinop = {({({(~WaitOnInput_inner_ready)}||(process_input[32]))}&&process_valid)}; 
  wire [64:0] WaitOnInput_inner_process_output;
  assign process_output = {{((WaitOnInput_inner_process_output[64])&&unnamedbinop36316USEDMULTIPLEbinop)},(WaitOnInput_inner_process_output[63:0])};
  // function: ready pure=true delay=0
  // function: reset pure=false delay=0
  // function: process pure=false delay=0
  ChangeRate_uint8_4_1__from1_to2_H1 #(.INSTANCE_NAME({INSTANCE_NAME,"_WaitOnInput_inner"})) WaitOnInput_inner(.CLK(CLK), .ready(WaitOnInput_inner_ready), .reset(reset), .CE(CE), .process_valid(unnamedbinop36316USEDMULTIPLEbinop), .process_input((process_input[31:0])), .process_output(WaitOnInput_inner_process_output));
endmodule

module LiftHandshake_WaitOnInput_ChangeRate_uint8_4_1__from1_to2_H1(input CLK, input ready_downstream, output ready, input reset, input [32:0] process_input, output [64:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire inner_WaitOnInput_ChangeRate_uint8_4_1__from1_to2_H1_ready;
  assign ready = {(inner_WaitOnInput_ChangeRate_uint8_4_1__from1_to2_H1_ready&&ready_downstream)};
  wire unnamedbinop36350USEDMULTIPLEbinop;assign unnamedbinop36350USEDMULTIPLEbinop = {(reset||ready_downstream)}; 
  wire unnamedunary36351USEDMULTIPLEunary;assign unnamedunary36351USEDMULTIPLEunary = {(~reset)}; 
  wire [64:0] inner_WaitOnInput_ChangeRate_uint8_4_1__from1_to2_H1_process_output;
  wire validBitDelay_WaitOnInput_ChangeRate_uint8_4_1__from1_to2_H1_pushPop_out;
  wire [64:0] unnamedtuple36361USEDMULTIPLEtuple;assign unnamedtuple36361USEDMULTIPLEtuple = {{((inner_WaitOnInput_ChangeRate_uint8_4_1__from1_to2_H1_process_output[64])&&validBitDelay_WaitOnInput_ChangeRate_uint8_4_1__from1_to2_H1_pushPop_out)},(inner_WaitOnInput_ChangeRate_uint8_4_1__from1_to2_H1_process_output[63:0])}; 
  always @(posedge CLK) begin if({(~{((unnamedtuple36361USEDMULTIPLEtuple[64])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: output valid bit should not be X!",INSTANCE_NAME); end end
  always @(posedge CLK) begin if({(~{((process_input[32])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = unnamedtuple36361USEDMULTIPLEtuple;
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  WaitOnInput_ChangeRate_uint8_4_1__from1_to2_H1 #(.INSTANCE_NAME({INSTANCE_NAME,"_inner_WaitOnInput_ChangeRate_uint8_4_1__from1_to2_H1"})) inner_WaitOnInput_ChangeRate_uint8_4_1__from1_to2_H1(.CLK(CLK), .ready(inner_WaitOnInput_ChangeRate_uint8_4_1__from1_to2_H1_ready), .reset(reset), .CE(unnamedbinop36350USEDMULTIPLEbinop), .process_valid(unnamedunary36351USEDMULTIPLEunary), .process_input(process_input), .process_output(inner_WaitOnInput_ChangeRate_uint8_4_1__from1_to2_H1_process_output));
  ShiftRegister_0_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_validBitDelay_WaitOnInput_ChangeRate_uint8_4_1__from1_to2_H1"})) validBitDelay_WaitOnInput_ChangeRate_uint8_4_1__from1_to2_H1(.CLK(CLK), .CE(unnamedbinop36350USEDMULTIPLEbinop), .sr_input((1'd1)), .pushPop_out(validBitDelay_WaitOnInput_ChangeRate_uint8_4_1__from1_to2_H1_pushPop_out));
endmodule

module sumwrap_uint16_to3(input CLK, input CE, input [31:0] process_input, output [15:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] unnamedcast49USEDMULTIPLEcast;assign unnamedcast49USEDMULTIPLEcast = (process_input[15:0]); 
  assign process_output = (({(unnamedcast49USEDMULTIPLEcast==(16'd3))})?((16'd0)):({(unnamedcast49USEDMULTIPLEcast+(process_input[31:16]))}));
  // function: process pure=true delay=0
endmodule

module RegBy_sumwrap_uint16_to3_CEtrue_initnil(input CLK, input set_valid, input CE, input [15:0] set_inp, input setby_valid, input [15:0] setby_inp, output [15:0] SETBY_OUTPUT, output [15:0] GET_OUTPUT);
parameter INSTANCE_NAME="INST";
  reg [15:0] R;
  wire [15:0] regby_inner_process_output;
  always @(posedge CLK) begin if(set_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(setby_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,set_valid})+({4'b0,setby_valid})) > 5'd1) begin $display("error, function 'set' on instance 'R' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [16:0] unnamedcallArbitrate89USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate89USEDMULTIPLEcallArbitrate = {(set_valid||setby_valid),((set_valid)?(set_inp):(regby_inner_process_output))}; 
    always @ (posedge CLK) begin if ((unnamedcallArbitrate89USEDMULTIPLEcallArbitrate[16]) && CE) begin R <= (unnamedcallArbitrate89USEDMULTIPLEcallArbitrate[15:0]); end end
  assign SETBY_OUTPUT = regby_inner_process_output;
  assign GET_OUTPUT = R;
  // function: set pure=false ONLY WIRE
  // function: setby pure=false ONLY WIRE
  // function: get pure=true ONLY WIRE
  sumwrap_uint16_to3 #(.INSTANCE_NAME({INSTANCE_NAME,"_regby_inner"})) regby_inner(.CLK(CLK), .CE(CE), .process_input({setby_inp,R}), .process_output(regby_inner_process_output));
endmodule

module ChangeRate_uint8_2_1__from4_to1_H1(input CLK, output ready, input reset, input CE, input process_valid, input [63:0] process_input, output [16:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  wire [15:0] phase_GET_OUTPUT;
  wire unnamedbinop100_readingUSEDMULTIPLEbinop;assign unnamedbinop100_readingUSEDMULTIPLEbinop = {(phase_GET_OUTPUT==(16'd0))}; 
  assign ready = unnamedbinop100_readingUSEDMULTIPLEbinop;
  reg [15:0] SR_2;
  wire [15:0] unnamedselect116USEDMULTIPLEselect;assign unnamedselect116USEDMULTIPLEselect = ((unnamedbinop100_readingUSEDMULTIPLEbinop)?(({process_input[15:0]})):(SR_2)); 
  reg [15:0] unnamedselect116_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect116_delay1_validunnamednull0_CECE <= unnamedselect116USEDMULTIPLEselect; end end
  reg [15:0] SR_1;  always @ (posedge CLK) begin if (process_valid && CE) begin SR_1 <= unnamedselect116USEDMULTIPLEselect; end end
  reg [15:0] SR_3;
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_2 <= ((unnamedbinop100_readingUSEDMULTIPLEbinop)?(({process_input[31:16]})):(SR_3)); end end
  reg [15:0] SR_4;
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_3 <= ((unnamedbinop100_readingUSEDMULTIPLEbinop)?(({process_input[47:32]})):(SR_4)); end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_4 <= ((unnamedbinop100_readingUSEDMULTIPLEbinop)?(({process_input[63:48]})):(SR_1)); end end
  wire [15:0] phase_SETBY_OUTPUT;
  assign process_output = {(1'd1),unnamedselect116_delay1_validunnamednull0_CECE};
  // function: ready pure=true delay=0
  // function: reset pure=false delay=0
  // function: process pure=false delay=1
  RegBy_sumwrap_uint16_to3_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_phase"})) phase(.CLK(CLK), .set_valid(reset), .CE(CE), .set_inp((16'd0)), .setby_valid(process_valid), .setby_inp((16'd1)), .SETBY_OUTPUT(phase_SETBY_OUTPUT), .GET_OUTPUT(phase_GET_OUTPUT));
endmodule

module WaitOnInput_ChangeRate_uint8_2_1__from4_to1_H1(input CLK, output ready, input reset, input CE, input process_valid, input [64:0] process_input, output [16:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  wire WaitOnInput_inner_ready;
  assign ready = WaitOnInput_inner_ready;
  wire unnamedbinop222USEDMULTIPLEbinop;assign unnamedbinop222USEDMULTIPLEbinop = {({({(~WaitOnInput_inner_ready)}||(process_input[64]))}&&process_valid)}; 
  wire [16:0] WaitOnInput_inner_process_output;
  reg unnamedbinop222_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedbinop222_delay1_validunnamednull0_CECE <= unnamedbinop222USEDMULTIPLEbinop; end end
  assign process_output = {{((WaitOnInput_inner_process_output[16])&&unnamedbinop222_delay1_validunnamednull0_CECE)},(WaitOnInput_inner_process_output[15:0])};
  // function: ready pure=true delay=0
  // function: reset pure=false delay=0
  // function: process pure=false delay=1
  ChangeRate_uint8_2_1__from4_to1_H1 #(.INSTANCE_NAME({INSTANCE_NAME,"_WaitOnInput_inner"})) WaitOnInput_inner(.CLK(CLK), .ready(WaitOnInput_inner_ready), .reset(reset), .CE(CE), .process_valid(unnamedbinop222USEDMULTIPLEbinop), .process_input((process_input[63:0])), .process_output(WaitOnInput_inner_process_output));
endmodule

module LiftHandshake_WaitOnInput_ChangeRate_uint8_2_1__from4_to1_H1(input CLK, input ready_downstream, output ready, input reset, input [64:0] process_input, output [16:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire inner_WaitOnInput_ChangeRate_uint8_2_1__from4_to1_H1_ready;
  assign ready = {(inner_WaitOnInput_ChangeRate_uint8_2_1__from4_to1_H1_ready&&ready_downstream)};
  wire unnamedbinop257USEDMULTIPLEbinop;assign unnamedbinop257USEDMULTIPLEbinop = {(reset||ready_downstream)}; 
  wire unnamedunary258USEDMULTIPLEunary;assign unnamedunary258USEDMULTIPLEunary = {(~reset)}; 
  wire [16:0] inner_WaitOnInput_ChangeRate_uint8_2_1__from4_to1_H1_process_output;
  wire validBitDelay_WaitOnInput_ChangeRate_uint8_2_1__from4_to1_H1_pushPop_out;
  wire [16:0] unnamedtuple290USEDMULTIPLEtuple;assign unnamedtuple290USEDMULTIPLEtuple = {{((inner_WaitOnInput_ChangeRate_uint8_2_1__from4_to1_H1_process_output[16])&&validBitDelay_WaitOnInput_ChangeRate_uint8_2_1__from4_to1_H1_pushPop_out)},(inner_WaitOnInput_ChangeRate_uint8_2_1__from4_to1_H1_process_output[15:0])}; 
  always @(posedge CLK) begin if({(~{((unnamedtuple290USEDMULTIPLEtuple[16])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: output valid bit should not be X!",INSTANCE_NAME); end end
  always @(posedge CLK) begin if({(~{((process_input[64])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = unnamedtuple290USEDMULTIPLEtuple;
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  WaitOnInput_ChangeRate_uint8_2_1__from4_to1_H1 #(.INSTANCE_NAME({INSTANCE_NAME,"_inner_WaitOnInput_ChangeRate_uint8_2_1__from4_to1_H1"})) inner_WaitOnInput_ChangeRate_uint8_2_1__from4_to1_H1(.CLK(CLK), .ready(inner_WaitOnInput_ChangeRate_uint8_2_1__from4_to1_H1_ready), .reset(reset), .CE(unnamedbinop257USEDMULTIPLEbinop), .process_valid(unnamedunary258USEDMULTIPLEunary), .process_input(process_input), .process_output(inner_WaitOnInput_ChangeRate_uint8_2_1__from4_to1_H1_process_output));
  ShiftRegister_1_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_validBitDelay_WaitOnInput_ChangeRate_uint8_2_1__from4_to1_H1"})) validBitDelay_WaitOnInput_ChangeRate_uint8_2_1__from4_to1_H1(.CLK(CLK), .pushPop_valid(unnamedunary258USEDMULTIPLEunary), .CE(unnamedbinop257USEDMULTIPLEbinop), .sr_input((1'd1)), .pushPop_out(validBitDelay_WaitOnInput_ChangeRate_uint8_2_1__from4_to1_H1_pushPop_out), .reset(reset));
endmodule

module PadSeq_uint8_2_1__W640_H480_L191_R0_B7_Top8_T11(input CLK, output ready, input reset, input CE, input process_valid, input [15:0] process_input, output [16:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  wire [15:0] posX_padSeq_GET_OUTPUT;
  wire [15:0] posY_padSeq_GET_OUTPUT;
  wire unnamedbinop441USEDMULTIPLEbinop;assign unnamedbinop441USEDMULTIPLEbinop = {({({((posX_padSeq_GET_OUTPUT)>=((16'd191)))}&&{((posX_padSeq_GET_OUTPUT)<((16'd831)))})}&&{({((posY_padSeq_GET_OUTPUT)>=((16'd7)))}&&{((posY_padSeq_GET_OUTPUT)<((16'd487)))})})}; 
  assign ready = unnamedbinop441USEDMULTIPLEbinop;
  reg [15:0] unnamedselect453_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect453_delay1_validunnamednull0_CECE <= ((unnamedbinop441USEDMULTIPLEbinop)?(process_input):({({8'd0, 8'd0})})); end end
  wire [15:0] posY_padSeq_SETBY_OUTPUT;
  wire [15:0] posX_padSeq_SETBY_OUTPUT;
  assign process_output = {(1'd1),unnamedselect453_delay1_validunnamednull0_CECE};
  // function: ready pure=true delay=0
  // function: reset pure=false delay=0
  // function: process pure=false delay=1
  RegBy_incif_wrapuint16_830_inc1_CEtrue_init0 #(.INSTANCE_NAME({INSTANCE_NAME,"_posX_padSeq"})) posX_padSeq(.CLK(CLK), .set_valid(reset), .CE(CE), .set_inp((16'd0)), .setby_valid(process_valid), .setby_inp((1'd1)), .SETBY_OUTPUT(posX_padSeq_SETBY_OUTPUT), .GET_OUTPUT(posX_padSeq_GET_OUTPUT));
  RegBy_incif_wrapuint16_494_incnil_CEtrue_init0 #(.INSTANCE_NAME({INSTANCE_NAME,"_posY_padSeq"})) posY_padSeq(.CLK(CLK), .set_valid(reset), .CE(CE), .set_inp((16'd0)), .setby_valid(process_valid), .setby_inp({(posX_padSeq_GET_OUTPUT==(16'd830))}), .SETBY_OUTPUT(posY_padSeq_SETBY_OUTPUT), .GET_OUTPUT(posY_padSeq_GET_OUTPUT));
endmodule

module WaitOnInput_PadSeq_uint8_2_1__W640_H480_L191_R0_B7_Top8_T11(input CLK, output ready, input reset, input CE, input process_valid, input [16:0] process_input, output [16:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  wire WaitOnInput_inner_ready;
  assign ready = WaitOnInput_inner_ready;
  wire unnamedbinop554USEDMULTIPLEbinop;assign unnamedbinop554USEDMULTIPLEbinop = {({({(~WaitOnInput_inner_ready)}||(process_input[16]))}&&process_valid)}; 
  wire [16:0] WaitOnInput_inner_process_output;
  reg unnamedbinop554_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedbinop554_delay1_validunnamednull0_CECE <= unnamedbinop554USEDMULTIPLEbinop; end end
  assign process_output = {{((WaitOnInput_inner_process_output[16])&&unnamedbinop554_delay1_validunnamednull0_CECE)},(WaitOnInput_inner_process_output[15:0])};
  // function: ready pure=true delay=0
  // function: reset pure=false delay=0
  // function: process pure=false delay=1
  PadSeq_uint8_2_1__W640_H480_L191_R0_B7_Top8_T11 #(.INSTANCE_NAME({INSTANCE_NAME,"_WaitOnInput_inner"})) WaitOnInput_inner(.CLK(CLK), .ready(WaitOnInput_inner_ready), .reset(reset), .CE(CE), .process_valid(unnamedbinop554USEDMULTIPLEbinop), .process_input((process_input[15:0])), .process_output(WaitOnInput_inner_process_output));
endmodule

module LiftHandshake_WaitOnInput_PadSeq_uint8_2_1__W640_H480_L191_R0_B7_Top8_T11(input CLK, input ready_downstream, output ready, input reset, input [16:0] process_input, output [16:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire inner_WaitOnInput_PadSeq_uint8_2_1__W640_H480_L191_R0_B7_Top8_T11_ready;
  assign ready = {(inner_WaitOnInput_PadSeq_uint8_2_1__W640_H480_L191_R0_B7_Top8_T11_ready&&ready_downstream)};
  wire unnamedbinop589USEDMULTIPLEbinop;assign unnamedbinop589USEDMULTIPLEbinop = {(reset||ready_downstream)}; 
  wire unnamedunary590USEDMULTIPLEunary;assign unnamedunary590USEDMULTIPLEunary = {(~reset)}; 
  wire [16:0] inner_WaitOnInput_PadSeq_uint8_2_1__W640_H480_L191_R0_B7_Top8_T11_process_output;
  wire validBitDelay_WaitOnInput_PadSeq_uint8_2_1__W640_H480_L191_R0_B7_Top8_T11_pushPop_out;
  wire [16:0] unnamedtuple600USEDMULTIPLEtuple;assign unnamedtuple600USEDMULTIPLEtuple = {{((inner_WaitOnInput_PadSeq_uint8_2_1__W640_H480_L191_R0_B7_Top8_T11_process_output[16])&&validBitDelay_WaitOnInput_PadSeq_uint8_2_1__W640_H480_L191_R0_B7_Top8_T11_pushPop_out)},(inner_WaitOnInput_PadSeq_uint8_2_1__W640_H480_L191_R0_B7_Top8_T11_process_output[15:0])}; 
  always @(posedge CLK) begin if({(~{((unnamedtuple600USEDMULTIPLEtuple[16])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: output valid bit should not be X!",INSTANCE_NAME); end end
  always @(posedge CLK) begin if({(~{((process_input[16])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = unnamedtuple600USEDMULTIPLEtuple;
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  WaitOnInput_PadSeq_uint8_2_1__W640_H480_L191_R0_B7_Top8_T11 #(.INSTANCE_NAME({INSTANCE_NAME,"_inner_WaitOnInput_PadSeq_uint8_2_1__W640_H480_L191_R0_B7_Top8_T11"})) inner_WaitOnInput_PadSeq_uint8_2_1__W640_H480_L191_R0_B7_Top8_T11(.CLK(CLK), .ready(inner_WaitOnInput_PadSeq_uint8_2_1__W640_H480_L191_R0_B7_Top8_T11_ready), .reset(reset), .CE(unnamedbinop589USEDMULTIPLEbinop), .process_valid(unnamedunary590USEDMULTIPLEunary), .process_input(process_input), .process_output(inner_WaitOnInput_PadSeq_uint8_2_1__W640_H480_L191_R0_B7_Top8_T11_process_output));
  ShiftRegister_1_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_validBitDelay_WaitOnInput_PadSeq_uint8_2_1__W640_H480_L191_R0_B7_Top8_T11"})) validBitDelay_WaitOnInput_PadSeq_uint8_2_1__W640_H480_L191_R0_B7_Top8_T11(.CLK(CLK), .pushPop_valid(unnamedunary590USEDMULTIPLEunary), .CE(unnamedbinop589USEDMULTIPLEbinop), .sr_input((1'd1)), .pushPop_out(validBitDelay_WaitOnInput_PadSeq_uint8_2_1__W640_H480_L191_R0_B7_Top8_T11_pushPop_out), .reset(reset));
endmodule

module slice_typeuint8_2_1__1_1__xl0_xh0_yl0_yh0(input CLK, input process_CE, input [15:0] inp, output [15:0] process_output);
parameter INSTANCE_NAME="INST";
  assign process_output = ({inp[15:0]});
  // function: process pure=true delay=0
endmodule

module MakeHandshake_slice_typeuint8_2_1__1_1__xl0_xh0_yl0_yh0(input CLK, input ready_downstream, output ready, input reset, input [16:0] process_input, output [16:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  assign ready = ready_downstream;
  wire unnamedbinop638USEDMULTIPLEbinop;assign unnamedbinop638USEDMULTIPLEbinop = {(ready_downstream||reset)}; 
  wire unnamedcast646USEDMULTIPLEcast;assign unnamedcast646USEDMULTIPLEcast = (process_input[16]); 
  wire [15:0] inner_process_output;
  wire validBitDelay_slice_typeuint8_2_1__1_1__xl0_xh0_yl0_yh0_pushPop_out;
  always @(posedge CLK) begin if({(~{(unnamedcast646USEDMULTIPLEcast===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: MakeHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = {validBitDelay_slice_typeuint8_2_1__1_1__xl0_xh0_yl0_yh0_pushPop_out,inner_process_output};
  // function: ready pure=true ONLY WIRE
  // function: reset pure=true ONLY WIRE
  // function: process pure=false ONLY WIRE
  ShiftRegister_0_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_validBitDelay_slice_typeuint8_2_1__1_1__xl0_xh0_yl0_yh0"})) validBitDelay_slice_typeuint8_2_1__1_1__xl0_xh0_yl0_yh0(.CLK(CLK), .CE(unnamedbinop638USEDMULTIPLEbinop), .sr_input(unnamedcast646USEDMULTIPLEcast), .pushPop_out(validBitDelay_slice_typeuint8_2_1__1_1__xl0_xh0_yl0_yh0_pushPop_out));
  slice_typeuint8_2_1__1_1__xl0_xh0_yl0_yh0 #(.INSTANCE_NAME({INSTANCE_NAME,"_inner"})) inner(.CLK(CLK), .process_CE(unnamedbinop638USEDMULTIPLEbinop), .inp((process_input[15:0])), .process_output(inner_process_output));
endmodule

module BroadcastStream_uint8_2_1__2(input CLK, input [1:0] ready_downstream, output ready, input reset_valid, input [16:0] process_input, output [33:0] process_output);
parameter INSTANCE_NAME="INST";
  wire unnamedbinop658USEDMULTIPLEbinop;assign unnamedbinop658USEDMULTIPLEbinop = {(({ready_downstream[0:0]})&&({ready_downstream[1:1]}))}; 
  assign ready = unnamedbinop658USEDMULTIPLEbinop;
  wire [16:0] unnamedtuple660USEDMULTIPLEtuple;assign unnamedtuple660USEDMULTIPLEtuple = {{((process_input[16])&&unnamedbinop658USEDMULTIPLEbinop)},(process_input[15:0])}; 
  assign process_output = {unnamedtuple660USEDMULTIPLEtuple,unnamedtuple660USEDMULTIPLEtuple};
  // function: ready pure=true ONLY WIRE
  // function: reset pure=true ONLY WIRE
  // function: process pure=true ONLY WIRE
endmodule

module slice_typeuint8_2_1__xl0_xh0_yl0_yh0(input CLK, input process_CE, input [15:0] inp, output [7:0] process_output);
parameter INSTANCE_NAME="INST";
  assign process_output = ({inp[7:0]});
  // function: process pure=true delay=0
endmodule

module MakeHandshake_slice_typeuint8_2_1__xl0_xh0_yl0_yh0(input CLK, input ready_downstream, output ready, input reset, input [16:0] process_input, output [8:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  assign ready = ready_downstream;
  wire unnamedbinop680USEDMULTIPLEbinop;assign unnamedbinop680USEDMULTIPLEbinop = {(ready_downstream||reset)}; 
  wire unnamedcast688USEDMULTIPLEcast;assign unnamedcast688USEDMULTIPLEcast = (process_input[16]); 
  wire [7:0] inner_process_output;
  wire validBitDelay_slice_typeuint8_2_1__xl0_xh0_yl0_yh0_pushPop_out;
  always @(posedge CLK) begin if({(~{(unnamedcast688USEDMULTIPLEcast===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: MakeHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = {validBitDelay_slice_typeuint8_2_1__xl0_xh0_yl0_yh0_pushPop_out,inner_process_output};
  // function: ready pure=true ONLY WIRE
  // function: reset pure=true ONLY WIRE
  // function: process pure=false ONLY WIRE
  ShiftRegister_0_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_validBitDelay_slice_typeuint8_2_1__xl0_xh0_yl0_yh0"})) validBitDelay_slice_typeuint8_2_1__xl0_xh0_yl0_yh0(.CLK(CLK), .CE(unnamedbinop680USEDMULTIPLEbinop), .sr_input(unnamedcast688USEDMULTIPLEcast), .pushPop_out(validBitDelay_slice_typeuint8_2_1__xl0_xh0_yl0_yh0_pushPop_out));
  slice_typeuint8_2_1__xl0_xh0_yl0_yh0 #(.INSTANCE_NAME({INSTANCE_NAME,"_inner"})) inner(.CLK(CLK), .process_CE(unnamedbinop680USEDMULTIPLEbinop), .inp((process_input[15:0])), .process_output(inner_process_output));
endmodule

module slice_typeuint8_2_1__xl1_xh1_yl0_yh0(input CLK, input process_CE, input [15:0] inp, output [7:0] process_output);
parameter INSTANCE_NAME="INST";
  assign process_output = ({inp[15:8]});
  // function: process pure=true delay=0
endmodule

module MakeHandshake_slice_typeuint8_2_1__xl1_xh1_yl0_yh0(input CLK, input ready_downstream, output ready, input reset, input [16:0] process_input, output [8:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  assign ready = ready_downstream;
  wire unnamedbinop21387USEDMULTIPLEbinop;assign unnamedbinop21387USEDMULTIPLEbinop = {(ready_downstream||reset)}; 
  wire unnamedcast21395USEDMULTIPLEcast;assign unnamedcast21395USEDMULTIPLEcast = (process_input[16]); 
  wire [7:0] inner_process_output;
  wire validBitDelay_slice_typeuint8_2_1__xl1_xh1_yl0_yh0_pushPop_out;
  always @(posedge CLK) begin if({(~{(unnamedcast21395USEDMULTIPLEcast===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: MakeHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = {validBitDelay_slice_typeuint8_2_1__xl1_xh1_yl0_yh0_pushPop_out,inner_process_output};
  // function: ready pure=true ONLY WIRE
  // function: reset pure=true ONLY WIRE
  // function: process pure=false ONLY WIRE
  ShiftRegister_0_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_validBitDelay_slice_typeuint8_2_1__xl1_xh1_yl0_yh0"})) validBitDelay_slice_typeuint8_2_1__xl1_xh1_yl0_yh0(.CLK(CLK), .CE(unnamedbinop21387USEDMULTIPLEbinop), .sr_input(unnamedcast21395USEDMULTIPLEcast), .pushPop_out(validBitDelay_slice_typeuint8_2_1__xl1_xh1_yl0_yh0_pushPop_out));
  slice_typeuint8_2_1__xl1_xh1_yl0_yh0 #(.INSTANCE_NAME({INSTANCE_NAME,"_inner"})) inner(.CLK(CLK), .process_CE(unnamedbinop21387USEDMULTIPLEbinop), .inp((process_input[15:0])), .process_output(inner_process_output));
endmodule

module arrayop_uint8_W1_Hnil(input CLK, input CE, input [7:0] process_input, output [7:0] process_output);
parameter INSTANCE_NAME="INST";
  assign process_output = {process_input};
  // function: process pure=true delay=0
  // function: reset pure=true delay=0
endmodule

module MakeHandshake_arrayop_uint8_W1_Hnil(input CLK, input ready_downstream, output ready, input reset, input [8:0] process_input, output [8:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  assign ready = ready_downstream;
  wire unnamedbinop1265USEDMULTIPLEbinop;assign unnamedbinop1265USEDMULTIPLEbinop = {(ready_downstream||reset)}; 
  wire unnamedcast1273USEDMULTIPLEcast;assign unnamedcast1273USEDMULTIPLEcast = (process_input[8]); 
  wire [7:0] inner_process_output;
  wire validBitDelay_arrayop_uint8_W1_Hnil_pushPop_out;
  always @(posedge CLK) begin if({(~{(unnamedcast1273USEDMULTIPLEcast===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: MakeHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = {validBitDelay_arrayop_uint8_W1_Hnil_pushPop_out,inner_process_output};
  // function: ready pure=true ONLY WIRE
  // function: reset pure=true ONLY WIRE
  // function: process pure=false ONLY WIRE
  ShiftRegister_0_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_validBitDelay_arrayop_uint8_W1_Hnil"})) validBitDelay_arrayop_uint8_W1_Hnil(.CLK(CLK), .CE(unnamedbinop1265USEDMULTIPLEbinop), .sr_input(unnamedcast1273USEDMULTIPLEcast), .pushPop_out(validBitDelay_arrayop_uint8_W1_Hnil_pushPop_out));
  arrayop_uint8_W1_Hnil #(.INSTANCE_NAME({INSTANCE_NAME,"_inner"})) inner(.CLK(CLK), .CE(unnamedbinop1265USEDMULTIPLEbinop), .process_input((process_input[7:0])), .process_output(inner_process_output));
endmodule

module ShiftRegister_15_CEtrue_TY1(input CLK, input pushPop_valid, input CE, input sr_input, output pushPop_out, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'pushPop'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  reg SR15;
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR1' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR1' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR1' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate2062USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate2062USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(sr_input):((1'd0)))}; 
  reg SR1;  always @ (posedge CLK) begin if ((unnamedcallArbitrate2062USEDMULTIPLEcallArbitrate[1]) && CE) begin SR1 <= (unnamedcallArbitrate2062USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR2' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR2' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR2' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate2068USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate2068USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR1):((1'd0)))}; 
  reg SR2;  always @ (posedge CLK) begin if ((unnamedcallArbitrate2068USEDMULTIPLEcallArbitrate[1]) && CE) begin SR2 <= (unnamedcallArbitrate2068USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR3' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR3' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR3' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate2074USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate2074USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR2):((1'd0)))}; 
  reg SR3;  always @ (posedge CLK) begin if ((unnamedcallArbitrate2074USEDMULTIPLEcallArbitrate[1]) && CE) begin SR3 <= (unnamedcallArbitrate2074USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR4' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR4' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR4' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate2080USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate2080USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR3):((1'd0)))}; 
  reg SR4;  always @ (posedge CLK) begin if ((unnamedcallArbitrate2080USEDMULTIPLEcallArbitrate[1]) && CE) begin SR4 <= (unnamedcallArbitrate2080USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR5' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR5' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR5' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate2086USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate2086USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR4):((1'd0)))}; 
  reg SR5;  always @ (posedge CLK) begin if ((unnamedcallArbitrate2086USEDMULTIPLEcallArbitrate[1]) && CE) begin SR5 <= (unnamedcallArbitrate2086USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR6' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR6' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR6' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate2092USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate2092USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR5):((1'd0)))}; 
  reg SR6;  always @ (posedge CLK) begin if ((unnamedcallArbitrate2092USEDMULTIPLEcallArbitrate[1]) && CE) begin SR6 <= (unnamedcallArbitrate2092USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR7' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR7' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR7' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate2098USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate2098USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR6):((1'd0)))}; 
  reg SR7;  always @ (posedge CLK) begin if ((unnamedcallArbitrate2098USEDMULTIPLEcallArbitrate[1]) && CE) begin SR7 <= (unnamedcallArbitrate2098USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR8' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR8' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR8' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate2104USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate2104USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR7):((1'd0)))}; 
  reg SR8;  always @ (posedge CLK) begin if ((unnamedcallArbitrate2104USEDMULTIPLEcallArbitrate[1]) && CE) begin SR8 <= (unnamedcallArbitrate2104USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR9' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR9' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR9' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate2110USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate2110USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR8):((1'd0)))}; 
  reg SR9;  always @ (posedge CLK) begin if ((unnamedcallArbitrate2110USEDMULTIPLEcallArbitrate[1]) && CE) begin SR9 <= (unnamedcallArbitrate2110USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR10' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR10' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR10' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate2116USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate2116USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR9):((1'd0)))}; 
  reg SR10;  always @ (posedge CLK) begin if ((unnamedcallArbitrate2116USEDMULTIPLEcallArbitrate[1]) && CE) begin SR10 <= (unnamedcallArbitrate2116USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR11' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR11' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR11' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate2122USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate2122USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR10):((1'd0)))}; 
  reg SR11;  always @ (posedge CLK) begin if ((unnamedcallArbitrate2122USEDMULTIPLEcallArbitrate[1]) && CE) begin SR11 <= (unnamedcallArbitrate2122USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR12' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR12' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR12' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate2128USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate2128USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR11):((1'd0)))}; 
  reg SR12;  always @ (posedge CLK) begin if ((unnamedcallArbitrate2128USEDMULTIPLEcallArbitrate[1]) && CE) begin SR12 <= (unnamedcallArbitrate2128USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR13' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR13' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR13' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate2134USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate2134USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR12):((1'd0)))}; 
  reg SR13;  always @ (posedge CLK) begin if ((unnamedcallArbitrate2134USEDMULTIPLEcallArbitrate[1]) && CE) begin SR13 <= (unnamedcallArbitrate2134USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR14' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR14' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR14' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate2140USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate2140USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR13):((1'd0)))}; 
  reg SR14;  always @ (posedge CLK) begin if ((unnamedcallArbitrate2140USEDMULTIPLEcallArbitrate[1]) && CE) begin SR14 <= (unnamedcallArbitrate2140USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR15' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR15' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR15' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate2146USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate2146USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR14):((1'd0)))}; 
    always @ (posedge CLK) begin if ((unnamedcallArbitrate2146USEDMULTIPLEcallArbitrate[1]) && CE) begin SR15 <= (unnamedcallArbitrate2146USEDMULTIPLEcallArbitrate[0]); end end
  assign pushPop_out = SR15;
  // function: pushPop pure=false delay=0
  // function: reset pure=false delay=0
endmodule

module incif_wrapuint16_830_incnil(input CLK, input CE, input [16:0] process_input, output [15:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] unnamedcast1278USEDMULTIPLEcast;assign unnamedcast1278USEDMULTIPLEcast = (process_input[15:0]); 
  assign process_output = (((process_input[16]))?((({(unnamedcast1278USEDMULTIPLEcast==(16'd830))})?((16'd0)):({(unnamedcast1278USEDMULTIPLEcast+(16'd1))}))):(unnamedcast1278USEDMULTIPLEcast));
  // function: process pure=true delay=0
endmodule

module RegBy_incif_wrapuint16_830_incnil_CEtrue_initnil(input CLK, input set_valid, input CE, input [15:0] set_inp, input setby_valid, input setby_inp, output [15:0] SETBY_OUTPUT, output [15:0] GET_OUTPUT);
parameter INSTANCE_NAME="INST";
  reg [15:0] R;
  wire [15:0] regby_inner_process_output;
  always @(posedge CLK) begin if(set_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(setby_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,set_valid})+({4'b0,setby_valid})) > 5'd1) begin $display("error, function 'set' on instance 'R' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [16:0] unnamedcallArbitrate1329USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate1329USEDMULTIPLEcallArbitrate = {(set_valid||setby_valid),((set_valid)?(set_inp):(regby_inner_process_output))}; 
    always @ (posedge CLK) begin if ((unnamedcallArbitrate1329USEDMULTIPLEcallArbitrate[16]) && CE) begin R <= (unnamedcallArbitrate1329USEDMULTIPLEcallArbitrate[15:0]); end end
  assign SETBY_OUTPUT = regby_inner_process_output;
  assign GET_OUTPUT = R;
  // function: set pure=false ONLY WIRE
  // function: setby pure=false ONLY WIRE
  // function: get pure=true ONLY WIRE
  incif_wrapuint16_830_incnil #(.INSTANCE_NAME({INSTANCE_NAME,"_regby_inner"})) regby_inner(.CLK(CLK), .CE(CE), .process_input({setby_inp,R}), .process_output(regby_inner_process_output));
endmodule

module bramSDP_WAROtrue_size1024_bw1_obwnil_CEtrue_initnil(input CLK, input writeAndReturnOriginal_valid, input writeAndReturnOriginal_CE, input [17:0] inp, output [7:0] WARO_OUT);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(writeAndReturnOriginal_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'writeAndReturnOriginal'", INSTANCE_NAME);  end end
  wire [7:0] unnamedcast1338;assign unnamedcast1338 = (inp[17:10]);  // wire for bitslice
  wire [7:0] bram_0_SET_AND_RETURN_ORIG_OUTPUT;
  assign WARO_OUT = {bram_0_SET_AND_RETURN_ORIG_OUTPUT};
  // function: writeAndReturnOriginal pure=false delay=1
  reg [7:0] bram_0_DI_B;
reg [10:0] bram_0_addr_B;
wire [7:0] bram_0_DO_B;
wire [18:0] bram_0_INPUT;
assign bram_0_INPUT = {unnamedcast1338[7:0],{1'b0,(inp[9:0])}};
RAMB16_S9_S9 #(.WRITE_MODE_A("READ_FIRST"),.WRITE_MODE_B("READ_FIRST")) bram_0 (
.DIPA(1'b0),
.DIPB(1'b0),
.DIA(bram_0_INPUT[18:11]),
.DIB(bram_0_DI_B),
.DOA(bram_0_SET_AND_RETURN_ORIG_OUTPUT),
.DOB(bram_0_DO_B),
.ADDRA(bram_0_INPUT[10:0]),
.ADDRB(bram_0_addr_B),
.WEA(writeAndReturnOriginal_valid),
.WEB(1'd0),
.ENA(writeAndReturnOriginal_CE),
.ENB(writeAndReturnOriginal_CE),
.CLKA(CLK),
.CLKB(CLK),
.SSRA(1'b0),
.SSRB(1'b0)
);


endmodule

module linebuffer_w831_h495_T1_ymin_15_Auint8(input CLK, input process_valid, input CE, input [7:0] process_input, output [127:0] process_output, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  wire [15:0] addr_GET_OUTPUT;
  wire [9:0] unnamedcast1506USEDMULTIPLEcast;assign unnamedcast1506USEDMULTIPLEcast = addr_GET_OUTPUT[9:0]; 
  reg [9:0] unnamedcast1506_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1506_delay1_validunnamednull0_CECE <= unnamedcast1506USEDMULTIPLEcast; end end
  reg [9:0] unnamedcast1506_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1506_delay2_validunnamednull0_CECE <= unnamedcast1506_delay1_validunnamednull0_CECE; end end
  reg [9:0] unnamedcast1506_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1506_delay3_validunnamednull0_CECE <= unnamedcast1506_delay2_validunnamednull0_CECE; end end
  reg [9:0] unnamedcast1506_delay4_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1506_delay4_validunnamednull0_CECE <= unnamedcast1506_delay3_validunnamednull0_CECE; end end
  reg [9:0] unnamedcast1506_delay5_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1506_delay5_validunnamednull0_CECE <= unnamedcast1506_delay4_validunnamednull0_CECE; end end
  reg [9:0] unnamedcast1506_delay6_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1506_delay6_validunnamednull0_CECE <= unnamedcast1506_delay5_validunnamednull0_CECE; end end
  reg [9:0] unnamedcast1506_delay7_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1506_delay7_validunnamednull0_CECE <= unnamedcast1506_delay6_validunnamednull0_CECE; end end
  reg [9:0] unnamedcast1506_delay8_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1506_delay8_validunnamednull0_CECE <= unnamedcast1506_delay7_validunnamednull0_CECE; end end
  reg [9:0] unnamedcast1506_delay9_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1506_delay9_validunnamednull0_CECE <= unnamedcast1506_delay8_validunnamednull0_CECE; end end
  reg [9:0] unnamedcast1506_delay10_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1506_delay10_validunnamednull0_CECE <= unnamedcast1506_delay9_validunnamednull0_CECE; end end
  reg [9:0] unnamedcast1506_delay11_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1506_delay11_validunnamednull0_CECE <= unnamedcast1506_delay10_validunnamednull0_CECE; end end
  reg [9:0] unnamedcast1506_delay12_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1506_delay12_validunnamednull0_CECE <= unnamedcast1506_delay11_validunnamednull0_CECE; end end
  reg [9:0] unnamedcast1506_delay13_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1506_delay13_validunnamednull0_CECE <= unnamedcast1506_delay12_validunnamednull0_CECE; end end
  reg [9:0] unnamedcast1506_delay14_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1506_delay14_validunnamednull0_CECE <= unnamedcast1506_delay13_validunnamednull0_CECE; end end
  wire [7:0] lb_m0_WARO_OUT;
  wire [7:0] unnamedcast1370USEDMULTIPLEcast;assign unnamedcast1370USEDMULTIPLEcast = lb_m0_WARO_OUT[7:0]; 
  reg process_valid_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay1_validunnamednull0_CECE <= process_valid; end end
  wire [7:0] lb_m1_WARO_OUT;
  wire [7:0] unnamedcast1380USEDMULTIPLEcast;assign unnamedcast1380USEDMULTIPLEcast = lb_m1_WARO_OUT[7:0]; 
  reg process_valid_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay2_validunnamednull0_CECE <= process_valid_delay1_validunnamednull0_CECE; end end
  wire [7:0] lb_m2_WARO_OUT;
  wire [7:0] unnamedcast1390USEDMULTIPLEcast;assign unnamedcast1390USEDMULTIPLEcast = lb_m2_WARO_OUT[7:0]; 
  reg process_valid_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay3_validunnamednull0_CECE <= process_valid_delay2_validunnamednull0_CECE; end end
  wire [7:0] lb_m3_WARO_OUT;
  wire [7:0] unnamedcast1400USEDMULTIPLEcast;assign unnamedcast1400USEDMULTIPLEcast = lb_m3_WARO_OUT[7:0]; 
  reg process_valid_delay4_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay4_validunnamednull0_CECE <= process_valid_delay3_validunnamednull0_CECE; end end
  wire [7:0] lb_m4_WARO_OUT;
  wire [7:0] unnamedcast1410USEDMULTIPLEcast;assign unnamedcast1410USEDMULTIPLEcast = lb_m4_WARO_OUT[7:0]; 
  reg process_valid_delay5_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay5_validunnamednull0_CECE <= process_valid_delay4_validunnamednull0_CECE; end end
  wire [7:0] lb_m5_WARO_OUT;
  wire [7:0] unnamedcast1420USEDMULTIPLEcast;assign unnamedcast1420USEDMULTIPLEcast = lb_m5_WARO_OUT[7:0]; 
  reg process_valid_delay6_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay6_validunnamednull0_CECE <= process_valid_delay5_validunnamednull0_CECE; end end
  wire [7:0] lb_m6_WARO_OUT;
  wire [7:0] unnamedcast1430USEDMULTIPLEcast;assign unnamedcast1430USEDMULTIPLEcast = lb_m6_WARO_OUT[7:0]; 
  reg process_valid_delay7_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay7_validunnamednull0_CECE <= process_valid_delay6_validunnamednull0_CECE; end end
  wire [7:0] lb_m7_WARO_OUT;
  wire [7:0] unnamedcast1440USEDMULTIPLEcast;assign unnamedcast1440USEDMULTIPLEcast = lb_m7_WARO_OUT[7:0]; 
  reg process_valid_delay8_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay8_validunnamednull0_CECE <= process_valid_delay7_validunnamednull0_CECE; end end
  wire [7:0] lb_m8_WARO_OUT;
  wire [7:0] unnamedcast1450USEDMULTIPLEcast;assign unnamedcast1450USEDMULTIPLEcast = lb_m8_WARO_OUT[7:0]; 
  reg process_valid_delay9_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay9_validunnamednull0_CECE <= process_valid_delay8_validunnamednull0_CECE; end end
  wire [7:0] lb_m9_WARO_OUT;
  wire [7:0] unnamedcast1460USEDMULTIPLEcast;assign unnamedcast1460USEDMULTIPLEcast = lb_m9_WARO_OUT[7:0]; 
  reg process_valid_delay10_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay10_validunnamednull0_CECE <= process_valid_delay9_validunnamednull0_CECE; end end
  wire [7:0] lb_m10_WARO_OUT;
  wire [7:0] unnamedcast1470USEDMULTIPLEcast;assign unnamedcast1470USEDMULTIPLEcast = lb_m10_WARO_OUT[7:0]; 
  reg process_valid_delay11_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay11_validunnamednull0_CECE <= process_valid_delay10_validunnamednull0_CECE; end end
  wire [7:0] lb_m11_WARO_OUT;
  wire [7:0] unnamedcast1480USEDMULTIPLEcast;assign unnamedcast1480USEDMULTIPLEcast = lb_m11_WARO_OUT[7:0]; 
  reg process_valid_delay12_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay12_validunnamednull0_CECE <= process_valid_delay11_validunnamednull0_CECE; end end
  wire [7:0] lb_m12_WARO_OUT;
  wire [7:0] unnamedcast1490USEDMULTIPLEcast;assign unnamedcast1490USEDMULTIPLEcast = lb_m12_WARO_OUT[7:0]; 
  reg process_valid_delay13_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay13_validunnamednull0_CECE <= process_valid_delay12_validunnamednull0_CECE; end end
  wire [7:0] lb_m13_WARO_OUT;
  wire [7:0] unnamedcast1500USEDMULTIPLEcast;assign unnamedcast1500USEDMULTIPLEcast = lb_m13_WARO_OUT[7:0]; 
  reg process_valid_delay14_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay14_validunnamednull0_CECE <= process_valid_delay13_validunnamednull0_CECE; end end
  wire [7:0] lb_m14_WARO_OUT;
  wire [7:0] unnamedcast1510;assign unnamedcast1510 = lb_m14_WARO_OUT[7:0];  // wire for array index
  reg [7:0] unnamedcast1502_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1502_delay1_validunnamednull0_CECE <= ({unnamedcast1500USEDMULTIPLEcast[7:0]}); end end
  reg [7:0] unnamedcast1492_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1492_delay1_validunnamednull0_CECE <= ({unnamedcast1490USEDMULTIPLEcast[7:0]}); end end
  reg [7:0] unnamedcast1492_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1492_delay2_validunnamednull0_CECE <= unnamedcast1492_delay1_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1482_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1482_delay1_validunnamednull0_CECE <= ({unnamedcast1480USEDMULTIPLEcast[7:0]}); end end
  reg [7:0] unnamedcast1482_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1482_delay2_validunnamednull0_CECE <= unnamedcast1482_delay1_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1482_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1482_delay3_validunnamednull0_CECE <= unnamedcast1482_delay2_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1472_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1472_delay1_validunnamednull0_CECE <= ({unnamedcast1470USEDMULTIPLEcast[7:0]}); end end
  reg [7:0] unnamedcast1472_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1472_delay2_validunnamednull0_CECE <= unnamedcast1472_delay1_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1472_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1472_delay3_validunnamednull0_CECE <= unnamedcast1472_delay2_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1472_delay4_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1472_delay4_validunnamednull0_CECE <= unnamedcast1472_delay3_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1462_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1462_delay1_validunnamednull0_CECE <= ({unnamedcast1460USEDMULTIPLEcast[7:0]}); end end
  reg [7:0] unnamedcast1462_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1462_delay2_validunnamednull0_CECE <= unnamedcast1462_delay1_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1462_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1462_delay3_validunnamednull0_CECE <= unnamedcast1462_delay2_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1462_delay4_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1462_delay4_validunnamednull0_CECE <= unnamedcast1462_delay3_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1462_delay5_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1462_delay5_validunnamednull0_CECE <= unnamedcast1462_delay4_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1452_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1452_delay1_validunnamednull0_CECE <= ({unnamedcast1450USEDMULTIPLEcast[7:0]}); end end
  reg [7:0] unnamedcast1452_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1452_delay2_validunnamednull0_CECE <= unnamedcast1452_delay1_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1452_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1452_delay3_validunnamednull0_CECE <= unnamedcast1452_delay2_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1452_delay4_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1452_delay4_validunnamednull0_CECE <= unnamedcast1452_delay3_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1452_delay5_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1452_delay5_validunnamednull0_CECE <= unnamedcast1452_delay4_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1452_delay6_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1452_delay6_validunnamednull0_CECE <= unnamedcast1452_delay5_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1442_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1442_delay1_validunnamednull0_CECE <= ({unnamedcast1440USEDMULTIPLEcast[7:0]}); end end
  reg [7:0] unnamedcast1442_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1442_delay2_validunnamednull0_CECE <= unnamedcast1442_delay1_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1442_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1442_delay3_validunnamednull0_CECE <= unnamedcast1442_delay2_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1442_delay4_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1442_delay4_validunnamednull0_CECE <= unnamedcast1442_delay3_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1442_delay5_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1442_delay5_validunnamednull0_CECE <= unnamedcast1442_delay4_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1442_delay6_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1442_delay6_validunnamednull0_CECE <= unnamedcast1442_delay5_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1442_delay7_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1442_delay7_validunnamednull0_CECE <= unnamedcast1442_delay6_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1432_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1432_delay1_validunnamednull0_CECE <= ({unnamedcast1430USEDMULTIPLEcast[7:0]}); end end
  reg [7:0] unnamedcast1432_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1432_delay2_validunnamednull0_CECE <= unnamedcast1432_delay1_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1432_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1432_delay3_validunnamednull0_CECE <= unnamedcast1432_delay2_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1432_delay4_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1432_delay4_validunnamednull0_CECE <= unnamedcast1432_delay3_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1432_delay5_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1432_delay5_validunnamednull0_CECE <= unnamedcast1432_delay4_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1432_delay6_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1432_delay6_validunnamednull0_CECE <= unnamedcast1432_delay5_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1432_delay7_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1432_delay7_validunnamednull0_CECE <= unnamedcast1432_delay6_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1432_delay8_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1432_delay8_validunnamednull0_CECE <= unnamedcast1432_delay7_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1422_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1422_delay1_validunnamednull0_CECE <= ({unnamedcast1420USEDMULTIPLEcast[7:0]}); end end
  reg [7:0] unnamedcast1422_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1422_delay2_validunnamednull0_CECE <= unnamedcast1422_delay1_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1422_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1422_delay3_validunnamednull0_CECE <= unnamedcast1422_delay2_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1422_delay4_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1422_delay4_validunnamednull0_CECE <= unnamedcast1422_delay3_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1422_delay5_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1422_delay5_validunnamednull0_CECE <= unnamedcast1422_delay4_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1422_delay6_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1422_delay6_validunnamednull0_CECE <= unnamedcast1422_delay5_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1422_delay7_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1422_delay7_validunnamednull0_CECE <= unnamedcast1422_delay6_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1422_delay8_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1422_delay8_validunnamednull0_CECE <= unnamedcast1422_delay7_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1422_delay9_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1422_delay9_validunnamednull0_CECE <= unnamedcast1422_delay8_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1412_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1412_delay1_validunnamednull0_CECE <= ({unnamedcast1410USEDMULTIPLEcast[7:0]}); end end
  reg [7:0] unnamedcast1412_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1412_delay2_validunnamednull0_CECE <= unnamedcast1412_delay1_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1412_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1412_delay3_validunnamednull0_CECE <= unnamedcast1412_delay2_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1412_delay4_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1412_delay4_validunnamednull0_CECE <= unnamedcast1412_delay3_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1412_delay5_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1412_delay5_validunnamednull0_CECE <= unnamedcast1412_delay4_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1412_delay6_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1412_delay6_validunnamednull0_CECE <= unnamedcast1412_delay5_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1412_delay7_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1412_delay7_validunnamednull0_CECE <= unnamedcast1412_delay6_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1412_delay8_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1412_delay8_validunnamednull0_CECE <= unnamedcast1412_delay7_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1412_delay9_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1412_delay9_validunnamednull0_CECE <= unnamedcast1412_delay8_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1412_delay10_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1412_delay10_validunnamednull0_CECE <= unnamedcast1412_delay9_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1402_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1402_delay1_validunnamednull0_CECE <= ({unnamedcast1400USEDMULTIPLEcast[7:0]}); end end
  reg [7:0] unnamedcast1402_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1402_delay2_validunnamednull0_CECE <= unnamedcast1402_delay1_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1402_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1402_delay3_validunnamednull0_CECE <= unnamedcast1402_delay2_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1402_delay4_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1402_delay4_validunnamednull0_CECE <= unnamedcast1402_delay3_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1402_delay5_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1402_delay5_validunnamednull0_CECE <= unnamedcast1402_delay4_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1402_delay6_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1402_delay6_validunnamednull0_CECE <= unnamedcast1402_delay5_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1402_delay7_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1402_delay7_validunnamednull0_CECE <= unnamedcast1402_delay6_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1402_delay8_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1402_delay8_validunnamednull0_CECE <= unnamedcast1402_delay7_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1402_delay9_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1402_delay9_validunnamednull0_CECE <= unnamedcast1402_delay8_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1402_delay10_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1402_delay10_validunnamednull0_CECE <= unnamedcast1402_delay9_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1402_delay11_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1402_delay11_validunnamednull0_CECE <= unnamedcast1402_delay10_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1392_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1392_delay1_validunnamednull0_CECE <= ({unnamedcast1390USEDMULTIPLEcast[7:0]}); end end
  reg [7:0] unnamedcast1392_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1392_delay2_validunnamednull0_CECE <= unnamedcast1392_delay1_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1392_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1392_delay3_validunnamednull0_CECE <= unnamedcast1392_delay2_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1392_delay4_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1392_delay4_validunnamednull0_CECE <= unnamedcast1392_delay3_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1392_delay5_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1392_delay5_validunnamednull0_CECE <= unnamedcast1392_delay4_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1392_delay6_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1392_delay6_validunnamednull0_CECE <= unnamedcast1392_delay5_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1392_delay7_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1392_delay7_validunnamednull0_CECE <= unnamedcast1392_delay6_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1392_delay8_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1392_delay8_validunnamednull0_CECE <= unnamedcast1392_delay7_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1392_delay9_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1392_delay9_validunnamednull0_CECE <= unnamedcast1392_delay8_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1392_delay10_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1392_delay10_validunnamednull0_CECE <= unnamedcast1392_delay9_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1392_delay11_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1392_delay11_validunnamednull0_CECE <= unnamedcast1392_delay10_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1392_delay12_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1392_delay12_validunnamednull0_CECE <= unnamedcast1392_delay11_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1382_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1382_delay1_validunnamednull0_CECE <= ({unnamedcast1380USEDMULTIPLEcast[7:0]}); end end
  reg [7:0] unnamedcast1382_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1382_delay2_validunnamednull0_CECE <= unnamedcast1382_delay1_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1382_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1382_delay3_validunnamednull0_CECE <= unnamedcast1382_delay2_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1382_delay4_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1382_delay4_validunnamednull0_CECE <= unnamedcast1382_delay3_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1382_delay5_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1382_delay5_validunnamednull0_CECE <= unnamedcast1382_delay4_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1382_delay6_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1382_delay6_validunnamednull0_CECE <= unnamedcast1382_delay5_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1382_delay7_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1382_delay7_validunnamednull0_CECE <= unnamedcast1382_delay6_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1382_delay8_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1382_delay8_validunnamednull0_CECE <= unnamedcast1382_delay7_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1382_delay9_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1382_delay9_validunnamednull0_CECE <= unnamedcast1382_delay8_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1382_delay10_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1382_delay10_validunnamednull0_CECE <= unnamedcast1382_delay9_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1382_delay11_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1382_delay11_validunnamednull0_CECE <= unnamedcast1382_delay10_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1382_delay12_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1382_delay12_validunnamednull0_CECE <= unnamedcast1382_delay11_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1382_delay13_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1382_delay13_validunnamednull0_CECE <= unnamedcast1382_delay12_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1372_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1372_delay1_validunnamednull0_CECE <= ({unnamedcast1370USEDMULTIPLEcast[7:0]}); end end
  reg [7:0] unnamedcast1372_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1372_delay2_validunnamednull0_CECE <= unnamedcast1372_delay1_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1372_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1372_delay3_validunnamednull0_CECE <= unnamedcast1372_delay2_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1372_delay4_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1372_delay4_validunnamednull0_CECE <= unnamedcast1372_delay3_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1372_delay5_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1372_delay5_validunnamednull0_CECE <= unnamedcast1372_delay4_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1372_delay6_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1372_delay6_validunnamednull0_CECE <= unnamedcast1372_delay5_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1372_delay7_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1372_delay7_validunnamednull0_CECE <= unnamedcast1372_delay6_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1372_delay8_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1372_delay8_validunnamednull0_CECE <= unnamedcast1372_delay7_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1372_delay9_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1372_delay9_validunnamednull0_CECE <= unnamedcast1372_delay8_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1372_delay10_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1372_delay10_validunnamednull0_CECE <= unnamedcast1372_delay9_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1372_delay11_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1372_delay11_validunnamednull0_CECE <= unnamedcast1372_delay10_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1372_delay12_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1372_delay12_validunnamednull0_CECE <= unnamedcast1372_delay11_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1372_delay13_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1372_delay13_validunnamednull0_CECE <= unnamedcast1372_delay12_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1372_delay14_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1372_delay14_validunnamednull0_CECE <= unnamedcast1372_delay13_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1346_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1346_delay1_validunnamednull0_CECE <= ({process_input[7:0]}); end end
  reg [7:0] unnamedcast1346_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1346_delay2_validunnamednull0_CECE <= unnamedcast1346_delay1_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1346_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1346_delay3_validunnamednull0_CECE <= unnamedcast1346_delay2_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1346_delay4_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1346_delay4_validunnamednull0_CECE <= unnamedcast1346_delay3_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1346_delay5_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1346_delay5_validunnamednull0_CECE <= unnamedcast1346_delay4_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1346_delay6_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1346_delay6_validunnamednull0_CECE <= unnamedcast1346_delay5_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1346_delay7_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1346_delay7_validunnamednull0_CECE <= unnamedcast1346_delay6_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1346_delay8_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1346_delay8_validunnamednull0_CECE <= unnamedcast1346_delay7_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1346_delay9_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1346_delay9_validunnamednull0_CECE <= unnamedcast1346_delay8_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1346_delay10_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1346_delay10_validunnamednull0_CECE <= unnamedcast1346_delay9_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1346_delay11_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1346_delay11_validunnamednull0_CECE <= unnamedcast1346_delay10_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1346_delay12_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1346_delay12_validunnamednull0_CECE <= unnamedcast1346_delay11_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1346_delay13_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1346_delay13_validunnamednull0_CECE <= unnamedcast1346_delay12_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1346_delay14_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1346_delay14_validunnamednull0_CECE <= unnamedcast1346_delay13_validunnamednull0_CECE; end end
  reg [7:0] unnamedcast1346_delay15_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast1346_delay15_validunnamednull0_CECE <= unnamedcast1346_delay14_validunnamednull0_CECE; end end
  wire [15:0] addr_SETBY_OUTPUT;
  assign process_output = {unnamedcast1346_delay15_validunnamednull0_CECE,unnamedcast1372_delay14_validunnamednull0_CECE,unnamedcast1382_delay13_validunnamednull0_CECE,unnamedcast1392_delay12_validunnamednull0_CECE,unnamedcast1402_delay11_validunnamednull0_CECE,unnamedcast1412_delay10_validunnamednull0_CECE,unnamedcast1422_delay9_validunnamednull0_CECE,unnamedcast1432_delay8_validunnamednull0_CECE,unnamedcast1442_delay7_validunnamednull0_CECE,unnamedcast1452_delay6_validunnamednull0_CECE,unnamedcast1462_delay5_validunnamednull0_CECE,unnamedcast1472_delay4_validunnamednull0_CECE,unnamedcast1482_delay3_validunnamednull0_CECE,unnamedcast1492_delay2_validunnamednull0_CECE,unnamedcast1502_delay1_validunnamednull0_CECE,({unnamedcast1510[7:0]})};
  // function: process pure=false delay=15
  // function: reset pure=false delay=0
  RegBy_incif_wrapuint16_830_incnil_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_addr"})) addr(.CLK(CLK), .set_valid(reset), .CE(CE), .set_inp((16'd0)), .setby_valid(process_valid), .setby_inp((1'd1)), .SETBY_OUTPUT(addr_SETBY_OUTPUT), .GET_OUTPUT(addr_GET_OUTPUT));
  bramSDP_WAROtrue_size1024_bw1_obwnil_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_lb_m0"})) lb_m0(.CLK(CLK), .writeAndReturnOriginal_valid(process_valid), .writeAndReturnOriginal_CE(CE), .inp({process_input,unnamedcast1506USEDMULTIPLEcast}), .WARO_OUT(lb_m0_WARO_OUT));
  bramSDP_WAROtrue_size1024_bw1_obwnil_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_lb_m1"})) lb_m1(.CLK(CLK), .writeAndReturnOriginal_valid(process_valid_delay1_validunnamednull0_CECE), .writeAndReturnOriginal_CE(CE), .inp({unnamedcast1370USEDMULTIPLEcast,unnamedcast1506_delay1_validunnamednull0_CECE}), .WARO_OUT(lb_m1_WARO_OUT));
  bramSDP_WAROtrue_size1024_bw1_obwnil_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_lb_m2"})) lb_m2(.CLK(CLK), .writeAndReturnOriginal_valid(process_valid_delay2_validunnamednull0_CECE), .writeAndReturnOriginal_CE(CE), .inp({unnamedcast1380USEDMULTIPLEcast,unnamedcast1506_delay2_validunnamednull0_CECE}), .WARO_OUT(lb_m2_WARO_OUT));
  bramSDP_WAROtrue_size1024_bw1_obwnil_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_lb_m3"})) lb_m3(.CLK(CLK), .writeAndReturnOriginal_valid(process_valid_delay3_validunnamednull0_CECE), .writeAndReturnOriginal_CE(CE), .inp({unnamedcast1390USEDMULTIPLEcast,unnamedcast1506_delay3_validunnamednull0_CECE}), .WARO_OUT(lb_m3_WARO_OUT));
  bramSDP_WAROtrue_size1024_bw1_obwnil_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_lb_m4"})) lb_m4(.CLK(CLK), .writeAndReturnOriginal_valid(process_valid_delay4_validunnamednull0_CECE), .writeAndReturnOriginal_CE(CE), .inp({unnamedcast1400USEDMULTIPLEcast,unnamedcast1506_delay4_validunnamednull0_CECE}), .WARO_OUT(lb_m4_WARO_OUT));
  bramSDP_WAROtrue_size1024_bw1_obwnil_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_lb_m5"})) lb_m5(.CLK(CLK), .writeAndReturnOriginal_valid(process_valid_delay5_validunnamednull0_CECE), .writeAndReturnOriginal_CE(CE), .inp({unnamedcast1410USEDMULTIPLEcast,unnamedcast1506_delay5_validunnamednull0_CECE}), .WARO_OUT(lb_m5_WARO_OUT));
  bramSDP_WAROtrue_size1024_bw1_obwnil_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_lb_m6"})) lb_m6(.CLK(CLK), .writeAndReturnOriginal_valid(process_valid_delay6_validunnamednull0_CECE), .writeAndReturnOriginal_CE(CE), .inp({unnamedcast1420USEDMULTIPLEcast,unnamedcast1506_delay6_validunnamednull0_CECE}), .WARO_OUT(lb_m6_WARO_OUT));
  bramSDP_WAROtrue_size1024_bw1_obwnil_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_lb_m7"})) lb_m7(.CLK(CLK), .writeAndReturnOriginal_valid(process_valid_delay7_validunnamednull0_CECE), .writeAndReturnOriginal_CE(CE), .inp({unnamedcast1430USEDMULTIPLEcast,unnamedcast1506_delay7_validunnamednull0_CECE}), .WARO_OUT(lb_m7_WARO_OUT));
  bramSDP_WAROtrue_size1024_bw1_obwnil_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_lb_m8"})) lb_m8(.CLK(CLK), .writeAndReturnOriginal_valid(process_valid_delay8_validunnamednull0_CECE), .writeAndReturnOriginal_CE(CE), .inp({unnamedcast1440USEDMULTIPLEcast,unnamedcast1506_delay8_validunnamednull0_CECE}), .WARO_OUT(lb_m8_WARO_OUT));
  bramSDP_WAROtrue_size1024_bw1_obwnil_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_lb_m9"})) lb_m9(.CLK(CLK), .writeAndReturnOriginal_valid(process_valid_delay9_validunnamednull0_CECE), .writeAndReturnOriginal_CE(CE), .inp({unnamedcast1450USEDMULTIPLEcast,unnamedcast1506_delay9_validunnamednull0_CECE}), .WARO_OUT(lb_m9_WARO_OUT));
  bramSDP_WAROtrue_size1024_bw1_obwnil_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_lb_m10"})) lb_m10(.CLK(CLK), .writeAndReturnOriginal_valid(process_valid_delay10_validunnamednull0_CECE), .writeAndReturnOriginal_CE(CE), .inp({unnamedcast1460USEDMULTIPLEcast,unnamedcast1506_delay10_validunnamednull0_CECE}), .WARO_OUT(lb_m10_WARO_OUT));
  bramSDP_WAROtrue_size1024_bw1_obwnil_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_lb_m11"})) lb_m11(.CLK(CLK), .writeAndReturnOriginal_valid(process_valid_delay11_validunnamednull0_CECE), .writeAndReturnOriginal_CE(CE), .inp({unnamedcast1470USEDMULTIPLEcast,unnamedcast1506_delay11_validunnamednull0_CECE}), .WARO_OUT(lb_m11_WARO_OUT));
  bramSDP_WAROtrue_size1024_bw1_obwnil_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_lb_m12"})) lb_m12(.CLK(CLK), .writeAndReturnOriginal_valid(process_valid_delay12_validunnamednull0_CECE), .writeAndReturnOriginal_CE(CE), .inp({unnamedcast1480USEDMULTIPLEcast,unnamedcast1506_delay12_validunnamednull0_CECE}), .WARO_OUT(lb_m12_WARO_OUT));
  bramSDP_WAROtrue_size1024_bw1_obwnil_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_lb_m13"})) lb_m13(.CLK(CLK), .writeAndReturnOriginal_valid(process_valid_delay13_validunnamednull0_CECE), .writeAndReturnOriginal_CE(CE), .inp({unnamedcast1490USEDMULTIPLEcast,unnamedcast1506_delay13_validunnamednull0_CECE}), .WARO_OUT(lb_m13_WARO_OUT));
  bramSDP_WAROtrue_size1024_bw1_obwnil_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_lb_m14"})) lb_m14(.CLK(CLK), .writeAndReturnOriginal_valid(process_valid_delay14_validunnamednull0_CECE), .writeAndReturnOriginal_CE(CE), .inp({unnamedcast1500USEDMULTIPLEcast,unnamedcast1506_delay14_validunnamednull0_CECE}), .WARO_OUT(lb_m14_WARO_OUT));
endmodule

module MakeHandshake_linebuffer_w831_h495_T1_ymin_15_Auint8(input CLK, input ready_downstream, output ready, input reset, input [8:0] process_input, output [128:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  assign ready = ready_downstream;
  wire unnamedbinop2158USEDMULTIPLEbinop;assign unnamedbinop2158USEDMULTIPLEbinop = {(ready_downstream||reset)}; 
  wire unnamedcast2166USEDMULTIPLEcast;assign unnamedcast2166USEDMULTIPLEcast = (process_input[8]); 
  wire [127:0] inner_process_output;
  wire validBitDelay_linebuffer_w831_h495_T1_ymin_15_Auint8_pushPop_out;
  always @(posedge CLK) begin if({(~{(unnamedcast2166USEDMULTIPLEcast===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: MakeHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = {validBitDelay_linebuffer_w831_h495_T1_ymin_15_Auint8_pushPop_out,inner_process_output};
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  ShiftRegister_15_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_validBitDelay_linebuffer_w831_h495_T1_ymin_15_Auint8"})) validBitDelay_linebuffer_w831_h495_T1_ymin_15_Auint8(.CLK(CLK), .pushPop_valid({(~reset)}), .CE(unnamedbinop2158USEDMULTIPLEbinop), .sr_input(unnamedcast2166USEDMULTIPLEcast), .pushPop_out(validBitDelay_linebuffer_w831_h495_T1_ymin_15_Auint8_pushPop_out), .reset(reset));
  linebuffer_w831_h495_T1_ymin_15_Auint8 #(.INSTANCE_NAME({INSTANCE_NAME,"_inner"})) inner(.CLK(CLK), .process_valid(unnamedcast2166USEDMULTIPLEcast), .CE(unnamedbinop2158USEDMULTIPLEbinop), .process_input((process_input[7:0])), .process_output(inner_process_output), .reset(reset));
endmodule

module sumwrap_uint16_to7(input CLK, input CE, input [31:0] process_input, output [15:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] unnamedcast2377USEDMULTIPLEcast;assign unnamedcast2377USEDMULTIPLEcast = (process_input[15:0]); 
  assign process_output = (({(unnamedcast2377USEDMULTIPLEcast==(16'd7))})?((16'd0)):({(unnamedcast2377USEDMULTIPLEcast+(process_input[31:16]))}));
  // function: process pure=true delay=0
endmodule

module RegBy_sumwrap_uint16_to7_CEtrue_initnil(input CLK, input set_valid, input CE, input [15:0] set_inp, input setby_valid, input [15:0] setby_inp, output [15:0] SETBY_OUTPUT, output [15:0] GET_OUTPUT);
parameter INSTANCE_NAME="INST";
  reg [15:0] R;
  wire [15:0] regby_inner_process_output;
  always @(posedge CLK) begin if(set_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(setby_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,set_valid})+({4'b0,setby_valid})) > 5'd1) begin $display("error, function 'set' on instance 'R' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [16:0] unnamedcallArbitrate2417USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate2417USEDMULTIPLEcallArbitrate = {(set_valid||setby_valid),((set_valid)?(set_inp):(regby_inner_process_output))}; 
    always @ (posedge CLK) begin if ((unnamedcallArbitrate2417USEDMULTIPLEcallArbitrate[16]) && CE) begin R <= (unnamedcallArbitrate2417USEDMULTIPLEcallArbitrate[15:0]); end end
  assign SETBY_OUTPUT = regby_inner_process_output;
  assign GET_OUTPUT = R;
  // function: set pure=false ONLY WIRE
  // function: setby pure=false ONLY WIRE
  // function: get pure=true ONLY WIRE
  sumwrap_uint16_to7 #(.INSTANCE_NAME({INSTANCE_NAME,"_regby_inner"})) regby_inner(.CLK(CLK), .CE(CE), .process_input({setby_inp,R}), .process_output(regby_inner_process_output));
endmodule

module SSRPartial_uint8_T0_125(input CLK, output ready, input reset, input CE, input process_valid, input [127:0] process_input, output [26368:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  wire [15:0] phase_GET_OUTPUT;
  wire unnamedbinop2428_readingUSEDMULTIPLEbinop;assign unnamedbinop2428_readingUSEDMULTIPLEbinop = {(phase_GET_OUTPUT==(16'd0))}; 
  assign ready = unnamedbinop2428_readingUSEDMULTIPLEbinop;
  reg [127:0] SR_194;
  reg [127:0] SR_3;
  wire [127:0] unnamedselect3255USEDMULTIPLEselect;assign unnamedselect3255USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_194):(SR_3)); 
  reg [127:0] unnamedselect3255_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3255_delay1_validunnamednull0_CECE <= unnamedselect3255USEDMULTIPLEselect; end end
  reg [127:0] SR_195;
  reg [127:0] SR_4;
  wire [127:0] unnamedselect3257USEDMULTIPLEselect;assign unnamedselect3257USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_195):(SR_4)); 
  reg [127:0] unnamedselect3257_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3257_delay1_validunnamednull0_CECE <= unnamedselect3257USEDMULTIPLEselect; end end
  reg [127:0] SR_196;
  reg [127:0] SR_5;
  wire [127:0] unnamedselect3259USEDMULTIPLEselect;assign unnamedselect3259USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_196):(SR_5)); 
  reg [127:0] unnamedselect3259_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3259_delay1_validunnamednull0_CECE <= unnamedselect3259USEDMULTIPLEselect; end end
  reg [127:0] SR_197;
  reg [127:0] SR_6;
  wire [127:0] unnamedselect3261USEDMULTIPLEselect;assign unnamedselect3261USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_197):(SR_6)); 
  reg [127:0] unnamedselect3261_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3261_delay1_validunnamednull0_CECE <= unnamedselect3261USEDMULTIPLEselect; end end
  reg [127:0] SR_198;
  reg [127:0] SR_7;
  wire [127:0] unnamedselect3263USEDMULTIPLEselect;assign unnamedselect3263USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_198):(SR_7)); 
  reg [127:0] unnamedselect3263_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3263_delay1_validunnamednull0_CECE <= unnamedselect3263USEDMULTIPLEselect; end end
  reg [127:0] SR_199;
  reg [127:0] SR_8;
  wire [127:0] unnamedselect3265USEDMULTIPLEselect;assign unnamedselect3265USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_199):(SR_8)); 
  reg [127:0] unnamedselect3265_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3265_delay1_validunnamednull0_CECE <= unnamedselect3265USEDMULTIPLEselect; end end
  reg [127:0] SR_200;
  reg [127:0] SR_9;
  wire [127:0] unnamedselect3267USEDMULTIPLEselect;assign unnamedselect3267USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_200):(SR_9)); 
  reg [127:0] unnamedselect3267_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3267_delay1_validunnamednull0_CECE <= unnamedselect3267USEDMULTIPLEselect; end end
  reg [127:0] SR_201;
  reg [127:0] SR_10;
  wire [127:0] unnamedselect3269USEDMULTIPLEselect;assign unnamedselect3269USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_201):(SR_10)); 
  reg [127:0] unnamedselect3269_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3269_delay1_validunnamednull0_CECE <= unnamedselect3269USEDMULTIPLEselect; end end
  reg [127:0] SR_202;
  reg [127:0] SR_11;
  wire [127:0] unnamedselect3271USEDMULTIPLEselect;assign unnamedselect3271USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_202):(SR_11)); 
  reg [127:0] unnamedselect3271_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3271_delay1_validunnamednull0_CECE <= unnamedselect3271USEDMULTIPLEselect; end end
  reg [127:0] SR_203;
  reg [127:0] SR_12;
  wire [127:0] unnamedselect3273USEDMULTIPLEselect;assign unnamedselect3273USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_203):(SR_12)); 
  reg [127:0] unnamedselect3273_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3273_delay1_validunnamednull0_CECE <= unnamedselect3273USEDMULTIPLEselect; end end
  reg [127:0] SR_204;
  reg [127:0] SR_13;
  wire [127:0] unnamedselect3275USEDMULTIPLEselect;assign unnamedselect3275USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_204):(SR_13)); 
  reg [127:0] unnamedselect3275_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3275_delay1_validunnamednull0_CECE <= unnamedselect3275USEDMULTIPLEselect; end end
  reg [127:0] SR_205;
  reg [127:0] SR_14;
  wire [127:0] unnamedselect3277USEDMULTIPLEselect;assign unnamedselect3277USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_205):(SR_14)); 
  reg [127:0] unnamedselect3277_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3277_delay1_validunnamednull0_CECE <= unnamedselect3277USEDMULTIPLEselect; end end
  reg [127:0] SR_206;
  reg [127:0] SR_15;
  wire [127:0] unnamedselect3279USEDMULTIPLEselect;assign unnamedselect3279USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_206):(SR_15)); 
  reg [127:0] unnamedselect3279_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3279_delay1_validunnamednull0_CECE <= unnamedselect3279USEDMULTIPLEselect; end end
  reg [127:0] SR_1;
  reg [127:0] SR_16;
  wire [127:0] unnamedselect3281USEDMULTIPLEselect;assign unnamedselect3281USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_1):(SR_16)); 
  reg [127:0] unnamedselect3281_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3281_delay1_validunnamednull0_CECE <= unnamedselect3281USEDMULTIPLEselect; end end
  reg [127:0] SR_2;
  reg [127:0] SR_17;
  wire [127:0] unnamedselect3283USEDMULTIPLEselect;assign unnamedselect3283USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_2):(SR_17)); 
  reg [127:0] unnamedselect3283_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3283_delay1_validunnamednull0_CECE <= unnamedselect3283USEDMULTIPLEselect; end end
  reg [127:0] SR_18;
  wire [127:0] unnamedselect3285USEDMULTIPLEselect;assign unnamedselect3285USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_3):(SR_18)); 
  reg [127:0] unnamedselect3285_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3285_delay1_validunnamednull0_CECE <= unnamedselect3285USEDMULTIPLEselect; end end
  reg [127:0] SR_19;
  wire [127:0] unnamedselect3287USEDMULTIPLEselect;assign unnamedselect3287USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_4):(SR_19)); 
  reg [127:0] unnamedselect3287_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3287_delay1_validunnamednull0_CECE <= unnamedselect3287USEDMULTIPLEselect; end end
  reg [127:0] SR_20;
  wire [127:0] unnamedselect3289USEDMULTIPLEselect;assign unnamedselect3289USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_5):(SR_20)); 
  reg [127:0] unnamedselect3289_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3289_delay1_validunnamednull0_CECE <= unnamedselect3289USEDMULTIPLEselect; end end
  reg [127:0] SR_21;
  wire [127:0] unnamedselect3291USEDMULTIPLEselect;assign unnamedselect3291USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_6):(SR_21)); 
  reg [127:0] unnamedselect3291_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3291_delay1_validunnamednull0_CECE <= unnamedselect3291USEDMULTIPLEselect; end end
  reg [127:0] SR_22;
  wire [127:0] unnamedselect3293USEDMULTIPLEselect;assign unnamedselect3293USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_7):(SR_22)); 
  reg [127:0] unnamedselect3293_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3293_delay1_validunnamednull0_CECE <= unnamedselect3293USEDMULTIPLEselect; end end
  reg [127:0] SR_23;
  wire [127:0] unnamedselect3295USEDMULTIPLEselect;assign unnamedselect3295USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_8):(SR_23)); 
  reg [127:0] unnamedselect3295_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3295_delay1_validunnamednull0_CECE <= unnamedselect3295USEDMULTIPLEselect; end end
  reg [127:0] SR_24;
  wire [127:0] unnamedselect3297USEDMULTIPLEselect;assign unnamedselect3297USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_9):(SR_24)); 
  reg [127:0] unnamedselect3297_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3297_delay1_validunnamednull0_CECE <= unnamedselect3297USEDMULTIPLEselect; end end
  reg [127:0] SR_25;
  wire [127:0] unnamedselect3299USEDMULTIPLEselect;assign unnamedselect3299USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_10):(SR_25)); 
  reg [127:0] unnamedselect3299_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3299_delay1_validunnamednull0_CECE <= unnamedselect3299USEDMULTIPLEselect; end end
  reg [127:0] SR_26;
  wire [127:0] unnamedselect3301USEDMULTIPLEselect;assign unnamedselect3301USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_11):(SR_26)); 
  reg [127:0] unnamedselect3301_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3301_delay1_validunnamednull0_CECE <= unnamedselect3301USEDMULTIPLEselect; end end
  reg [127:0] SR_27;
  wire [127:0] unnamedselect3303USEDMULTIPLEselect;assign unnamedselect3303USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_12):(SR_27)); 
  reg [127:0] unnamedselect3303_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3303_delay1_validunnamednull0_CECE <= unnamedselect3303USEDMULTIPLEselect; end end
  reg [127:0] SR_28;
  wire [127:0] unnamedselect3305USEDMULTIPLEselect;assign unnamedselect3305USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_13):(SR_28)); 
  reg [127:0] unnamedselect3305_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3305_delay1_validunnamednull0_CECE <= unnamedselect3305USEDMULTIPLEselect; end end
  reg [127:0] SR_29;
  wire [127:0] unnamedselect3307USEDMULTIPLEselect;assign unnamedselect3307USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_14):(SR_29)); 
  reg [127:0] unnamedselect3307_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3307_delay1_validunnamednull0_CECE <= unnamedselect3307USEDMULTIPLEselect; end end
  reg [127:0] SR_30;
  wire [127:0] unnamedselect3309USEDMULTIPLEselect;assign unnamedselect3309USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_15):(SR_30)); 
  reg [127:0] unnamedselect3309_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3309_delay1_validunnamednull0_CECE <= unnamedselect3309USEDMULTIPLEselect; end end
  reg [127:0] SR_31;
  wire [127:0] unnamedselect3311USEDMULTIPLEselect;assign unnamedselect3311USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_16):(SR_31)); 
  reg [127:0] unnamedselect3311_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3311_delay1_validunnamednull0_CECE <= unnamedselect3311USEDMULTIPLEselect; end end
  reg [127:0] SR_32;
  wire [127:0] unnamedselect3313USEDMULTIPLEselect;assign unnamedselect3313USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_17):(SR_32)); 
  reg [127:0] unnamedselect3313_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3313_delay1_validunnamednull0_CECE <= unnamedselect3313USEDMULTIPLEselect; end end
  reg [127:0] SR_33;
  wire [127:0] unnamedselect3315USEDMULTIPLEselect;assign unnamedselect3315USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_18):(SR_33)); 
  reg [127:0] unnamedselect3315_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3315_delay1_validunnamednull0_CECE <= unnamedselect3315USEDMULTIPLEselect; end end
  reg [127:0] SR_34;
  wire [127:0] unnamedselect3317USEDMULTIPLEselect;assign unnamedselect3317USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_19):(SR_34)); 
  reg [127:0] unnamedselect3317_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3317_delay1_validunnamednull0_CECE <= unnamedselect3317USEDMULTIPLEselect; end end
  reg [127:0] SR_35;
  wire [127:0] unnamedselect3319USEDMULTIPLEselect;assign unnamedselect3319USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_20):(SR_35)); 
  reg [127:0] unnamedselect3319_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3319_delay1_validunnamednull0_CECE <= unnamedselect3319USEDMULTIPLEselect; end end
  reg [127:0] SR_36;
  wire [127:0] unnamedselect3321USEDMULTIPLEselect;assign unnamedselect3321USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_21):(SR_36)); 
  reg [127:0] unnamedselect3321_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3321_delay1_validunnamednull0_CECE <= unnamedselect3321USEDMULTIPLEselect; end end
  reg [127:0] SR_37;
  wire [127:0] unnamedselect3323USEDMULTIPLEselect;assign unnamedselect3323USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_22):(SR_37)); 
  reg [127:0] unnamedselect3323_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3323_delay1_validunnamednull0_CECE <= unnamedselect3323USEDMULTIPLEselect; end end
  reg [127:0] SR_38;
  wire [127:0] unnamedselect3325USEDMULTIPLEselect;assign unnamedselect3325USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_23):(SR_38)); 
  reg [127:0] unnamedselect3325_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3325_delay1_validunnamednull0_CECE <= unnamedselect3325USEDMULTIPLEselect; end end
  reg [127:0] SR_39;
  wire [127:0] unnamedselect3327USEDMULTIPLEselect;assign unnamedselect3327USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_24):(SR_39)); 
  reg [127:0] unnamedselect3327_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3327_delay1_validunnamednull0_CECE <= unnamedselect3327USEDMULTIPLEselect; end end
  reg [127:0] SR_40;
  wire [127:0] unnamedselect3329USEDMULTIPLEselect;assign unnamedselect3329USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_25):(SR_40)); 
  reg [127:0] unnamedselect3329_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3329_delay1_validunnamednull0_CECE <= unnamedselect3329USEDMULTIPLEselect; end end
  reg [127:0] SR_41;
  wire [127:0] unnamedselect3331USEDMULTIPLEselect;assign unnamedselect3331USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_26):(SR_41)); 
  reg [127:0] unnamedselect3331_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3331_delay1_validunnamednull0_CECE <= unnamedselect3331USEDMULTIPLEselect; end end
  reg [127:0] SR_42;
  wire [127:0] unnamedselect3333USEDMULTIPLEselect;assign unnamedselect3333USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_27):(SR_42)); 
  reg [127:0] unnamedselect3333_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3333_delay1_validunnamednull0_CECE <= unnamedselect3333USEDMULTIPLEselect; end end
  reg [127:0] SR_43;
  wire [127:0] unnamedselect3335USEDMULTIPLEselect;assign unnamedselect3335USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_28):(SR_43)); 
  reg [127:0] unnamedselect3335_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3335_delay1_validunnamednull0_CECE <= unnamedselect3335USEDMULTIPLEselect; end end
  reg [127:0] SR_44;
  wire [127:0] unnamedselect3337USEDMULTIPLEselect;assign unnamedselect3337USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_29):(SR_44)); 
  reg [127:0] unnamedselect3337_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3337_delay1_validunnamednull0_CECE <= unnamedselect3337USEDMULTIPLEselect; end end
  reg [127:0] SR_45;
  wire [127:0] unnamedselect3339USEDMULTIPLEselect;assign unnamedselect3339USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_30):(SR_45)); 
  reg [127:0] unnamedselect3339_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3339_delay1_validunnamednull0_CECE <= unnamedselect3339USEDMULTIPLEselect; end end
  reg [127:0] SR_46;
  wire [127:0] unnamedselect3341USEDMULTIPLEselect;assign unnamedselect3341USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_31):(SR_46)); 
  reg [127:0] unnamedselect3341_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3341_delay1_validunnamednull0_CECE <= unnamedselect3341USEDMULTIPLEselect; end end
  reg [127:0] SR_47;
  wire [127:0] unnamedselect3343USEDMULTIPLEselect;assign unnamedselect3343USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_32):(SR_47)); 
  reg [127:0] unnamedselect3343_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3343_delay1_validunnamednull0_CECE <= unnamedselect3343USEDMULTIPLEselect; end end
  reg [127:0] SR_48;
  wire [127:0] unnamedselect3345USEDMULTIPLEselect;assign unnamedselect3345USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_33):(SR_48)); 
  reg [127:0] unnamedselect3345_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3345_delay1_validunnamednull0_CECE <= unnamedselect3345USEDMULTIPLEselect; end end
  reg [127:0] SR_49;
  wire [127:0] unnamedselect3347USEDMULTIPLEselect;assign unnamedselect3347USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_34):(SR_49)); 
  reg [127:0] unnamedselect3347_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3347_delay1_validunnamednull0_CECE <= unnamedselect3347USEDMULTIPLEselect; end end
  reg [127:0] SR_50;
  wire [127:0] unnamedselect3349USEDMULTIPLEselect;assign unnamedselect3349USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_35):(SR_50)); 
  reg [127:0] unnamedselect3349_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3349_delay1_validunnamednull0_CECE <= unnamedselect3349USEDMULTIPLEselect; end end
  reg [127:0] SR_51;
  wire [127:0] unnamedselect3351USEDMULTIPLEselect;assign unnamedselect3351USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_36):(SR_51)); 
  reg [127:0] unnamedselect3351_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3351_delay1_validunnamednull0_CECE <= unnamedselect3351USEDMULTIPLEselect; end end
  reg [127:0] SR_52;
  wire [127:0] unnamedselect3353USEDMULTIPLEselect;assign unnamedselect3353USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_37):(SR_52)); 
  reg [127:0] unnamedselect3353_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3353_delay1_validunnamednull0_CECE <= unnamedselect3353USEDMULTIPLEselect; end end
  reg [127:0] SR_53;
  wire [127:0] unnamedselect3355USEDMULTIPLEselect;assign unnamedselect3355USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_38):(SR_53)); 
  reg [127:0] unnamedselect3355_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3355_delay1_validunnamednull0_CECE <= unnamedselect3355USEDMULTIPLEselect; end end
  reg [127:0] SR_54;
  wire [127:0] unnamedselect3357USEDMULTIPLEselect;assign unnamedselect3357USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_39):(SR_54)); 
  reg [127:0] unnamedselect3357_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3357_delay1_validunnamednull0_CECE <= unnamedselect3357USEDMULTIPLEselect; end end
  reg [127:0] SR_55;
  wire [127:0] unnamedselect3359USEDMULTIPLEselect;assign unnamedselect3359USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_40):(SR_55)); 
  reg [127:0] unnamedselect3359_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3359_delay1_validunnamednull0_CECE <= unnamedselect3359USEDMULTIPLEselect; end end
  reg [127:0] SR_56;
  wire [127:0] unnamedselect3361USEDMULTIPLEselect;assign unnamedselect3361USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_41):(SR_56)); 
  reg [127:0] unnamedselect3361_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3361_delay1_validunnamednull0_CECE <= unnamedselect3361USEDMULTIPLEselect; end end
  reg [127:0] SR_57;
  wire [127:0] unnamedselect3363USEDMULTIPLEselect;assign unnamedselect3363USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_42):(SR_57)); 
  reg [127:0] unnamedselect3363_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3363_delay1_validunnamednull0_CECE <= unnamedselect3363USEDMULTIPLEselect; end end
  reg [127:0] SR_58;
  wire [127:0] unnamedselect3365USEDMULTIPLEselect;assign unnamedselect3365USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_43):(SR_58)); 
  reg [127:0] unnamedselect3365_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3365_delay1_validunnamednull0_CECE <= unnamedselect3365USEDMULTIPLEselect; end end
  reg [127:0] SR_59;
  wire [127:0] unnamedselect3367USEDMULTIPLEselect;assign unnamedselect3367USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_44):(SR_59)); 
  reg [127:0] unnamedselect3367_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3367_delay1_validunnamednull0_CECE <= unnamedselect3367USEDMULTIPLEselect; end end
  reg [127:0] SR_60;
  wire [127:0] unnamedselect3369USEDMULTIPLEselect;assign unnamedselect3369USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_45):(SR_60)); 
  reg [127:0] unnamedselect3369_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3369_delay1_validunnamednull0_CECE <= unnamedselect3369USEDMULTIPLEselect; end end
  reg [127:0] SR_61;
  wire [127:0] unnamedselect3371USEDMULTIPLEselect;assign unnamedselect3371USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_46):(SR_61)); 
  reg [127:0] unnamedselect3371_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3371_delay1_validunnamednull0_CECE <= unnamedselect3371USEDMULTIPLEselect; end end
  reg [127:0] SR_62;
  wire [127:0] unnamedselect3373USEDMULTIPLEselect;assign unnamedselect3373USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_47):(SR_62)); 
  reg [127:0] unnamedselect3373_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3373_delay1_validunnamednull0_CECE <= unnamedselect3373USEDMULTIPLEselect; end end
  reg [127:0] SR_63;
  wire [127:0] unnamedselect3375USEDMULTIPLEselect;assign unnamedselect3375USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_48):(SR_63)); 
  reg [127:0] unnamedselect3375_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3375_delay1_validunnamednull0_CECE <= unnamedselect3375USEDMULTIPLEselect; end end
  reg [127:0] SR_64;
  wire [127:0] unnamedselect3377USEDMULTIPLEselect;assign unnamedselect3377USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_49):(SR_64)); 
  reg [127:0] unnamedselect3377_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3377_delay1_validunnamednull0_CECE <= unnamedselect3377USEDMULTIPLEselect; end end
  reg [127:0] SR_65;
  wire [127:0] unnamedselect3379USEDMULTIPLEselect;assign unnamedselect3379USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_50):(SR_65)); 
  reg [127:0] unnamedselect3379_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3379_delay1_validunnamednull0_CECE <= unnamedselect3379USEDMULTIPLEselect; end end
  reg [127:0] SR_66;
  wire [127:0] unnamedselect3381USEDMULTIPLEselect;assign unnamedselect3381USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_51):(SR_66)); 
  reg [127:0] unnamedselect3381_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3381_delay1_validunnamednull0_CECE <= unnamedselect3381USEDMULTIPLEselect; end end
  reg [127:0] SR_67;
  wire [127:0] unnamedselect3383USEDMULTIPLEselect;assign unnamedselect3383USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_52):(SR_67)); 
  reg [127:0] unnamedselect3383_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3383_delay1_validunnamednull0_CECE <= unnamedselect3383USEDMULTIPLEselect; end end
  reg [127:0] SR_68;
  wire [127:0] unnamedselect3385USEDMULTIPLEselect;assign unnamedselect3385USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_53):(SR_68)); 
  reg [127:0] unnamedselect3385_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3385_delay1_validunnamednull0_CECE <= unnamedselect3385USEDMULTIPLEselect; end end
  reg [127:0] SR_69;
  wire [127:0] unnamedselect3387USEDMULTIPLEselect;assign unnamedselect3387USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_54):(SR_69)); 
  reg [127:0] unnamedselect3387_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3387_delay1_validunnamednull0_CECE <= unnamedselect3387USEDMULTIPLEselect; end end
  reg [127:0] SR_70;
  wire [127:0] unnamedselect3389USEDMULTIPLEselect;assign unnamedselect3389USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_55):(SR_70)); 
  reg [127:0] unnamedselect3389_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3389_delay1_validunnamednull0_CECE <= unnamedselect3389USEDMULTIPLEselect; end end
  reg [127:0] SR_71;
  wire [127:0] unnamedselect3391USEDMULTIPLEselect;assign unnamedselect3391USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_56):(SR_71)); 
  reg [127:0] unnamedselect3391_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3391_delay1_validunnamednull0_CECE <= unnamedselect3391USEDMULTIPLEselect; end end
  reg [127:0] SR_72;
  wire [127:0] unnamedselect3393USEDMULTIPLEselect;assign unnamedselect3393USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_57):(SR_72)); 
  reg [127:0] unnamedselect3393_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3393_delay1_validunnamednull0_CECE <= unnamedselect3393USEDMULTIPLEselect; end end
  reg [127:0] SR_73;
  wire [127:0] unnamedselect3395USEDMULTIPLEselect;assign unnamedselect3395USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_58):(SR_73)); 
  reg [127:0] unnamedselect3395_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3395_delay1_validunnamednull0_CECE <= unnamedselect3395USEDMULTIPLEselect; end end
  reg [127:0] SR_74;
  wire [127:0] unnamedselect3397USEDMULTIPLEselect;assign unnamedselect3397USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_59):(SR_74)); 
  reg [127:0] unnamedselect3397_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3397_delay1_validunnamednull0_CECE <= unnamedselect3397USEDMULTIPLEselect; end end
  reg [127:0] SR_75;
  wire [127:0] unnamedselect3399USEDMULTIPLEselect;assign unnamedselect3399USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_60):(SR_75)); 
  reg [127:0] unnamedselect3399_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3399_delay1_validunnamednull0_CECE <= unnamedselect3399USEDMULTIPLEselect; end end
  reg [127:0] SR_76;
  wire [127:0] unnamedselect3401USEDMULTIPLEselect;assign unnamedselect3401USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_61):(SR_76)); 
  reg [127:0] unnamedselect3401_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3401_delay1_validunnamednull0_CECE <= unnamedselect3401USEDMULTIPLEselect; end end
  reg [127:0] SR_77;
  wire [127:0] unnamedselect3403USEDMULTIPLEselect;assign unnamedselect3403USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_62):(SR_77)); 
  reg [127:0] unnamedselect3403_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3403_delay1_validunnamednull0_CECE <= unnamedselect3403USEDMULTIPLEselect; end end
  reg [127:0] SR_78;
  wire [127:0] unnamedselect3405USEDMULTIPLEselect;assign unnamedselect3405USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_63):(SR_78)); 
  reg [127:0] unnamedselect3405_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3405_delay1_validunnamednull0_CECE <= unnamedselect3405USEDMULTIPLEselect; end end
  reg [127:0] SR_79;
  wire [127:0] unnamedselect3407USEDMULTIPLEselect;assign unnamedselect3407USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_64):(SR_79)); 
  reg [127:0] unnamedselect3407_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3407_delay1_validunnamednull0_CECE <= unnamedselect3407USEDMULTIPLEselect; end end
  reg [127:0] SR_80;
  wire [127:0] unnamedselect3409USEDMULTIPLEselect;assign unnamedselect3409USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_65):(SR_80)); 
  reg [127:0] unnamedselect3409_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3409_delay1_validunnamednull0_CECE <= unnamedselect3409USEDMULTIPLEselect; end end
  reg [127:0] SR_81;
  wire [127:0] unnamedselect3411USEDMULTIPLEselect;assign unnamedselect3411USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_66):(SR_81)); 
  reg [127:0] unnamedselect3411_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3411_delay1_validunnamednull0_CECE <= unnamedselect3411USEDMULTIPLEselect; end end
  reg [127:0] SR_82;
  wire [127:0] unnamedselect3413USEDMULTIPLEselect;assign unnamedselect3413USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_67):(SR_82)); 
  reg [127:0] unnamedselect3413_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3413_delay1_validunnamednull0_CECE <= unnamedselect3413USEDMULTIPLEselect; end end
  reg [127:0] SR_83;
  wire [127:0] unnamedselect3415USEDMULTIPLEselect;assign unnamedselect3415USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_68):(SR_83)); 
  reg [127:0] unnamedselect3415_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3415_delay1_validunnamednull0_CECE <= unnamedselect3415USEDMULTIPLEselect; end end
  reg [127:0] SR_84;
  wire [127:0] unnamedselect3417USEDMULTIPLEselect;assign unnamedselect3417USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_69):(SR_84)); 
  reg [127:0] unnamedselect3417_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3417_delay1_validunnamednull0_CECE <= unnamedselect3417USEDMULTIPLEselect; end end
  reg [127:0] SR_85;
  wire [127:0] unnamedselect3419USEDMULTIPLEselect;assign unnamedselect3419USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_70):(SR_85)); 
  reg [127:0] unnamedselect3419_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3419_delay1_validunnamednull0_CECE <= unnamedselect3419USEDMULTIPLEselect; end end
  reg [127:0] SR_86;
  wire [127:0] unnamedselect3421USEDMULTIPLEselect;assign unnamedselect3421USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_71):(SR_86)); 
  reg [127:0] unnamedselect3421_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3421_delay1_validunnamednull0_CECE <= unnamedselect3421USEDMULTIPLEselect; end end
  reg [127:0] SR_87;
  wire [127:0] unnamedselect3423USEDMULTIPLEselect;assign unnamedselect3423USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_72):(SR_87)); 
  reg [127:0] unnamedselect3423_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3423_delay1_validunnamednull0_CECE <= unnamedselect3423USEDMULTIPLEselect; end end
  reg [127:0] SR_88;
  wire [127:0] unnamedselect3425USEDMULTIPLEselect;assign unnamedselect3425USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_73):(SR_88)); 
  reg [127:0] unnamedselect3425_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3425_delay1_validunnamednull0_CECE <= unnamedselect3425USEDMULTIPLEselect; end end
  reg [127:0] SR_89;
  wire [127:0] unnamedselect3427USEDMULTIPLEselect;assign unnamedselect3427USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_74):(SR_89)); 
  reg [127:0] unnamedselect3427_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3427_delay1_validunnamednull0_CECE <= unnamedselect3427USEDMULTIPLEselect; end end
  reg [127:0] SR_90;
  wire [127:0] unnamedselect3429USEDMULTIPLEselect;assign unnamedselect3429USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_75):(SR_90)); 
  reg [127:0] unnamedselect3429_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3429_delay1_validunnamednull0_CECE <= unnamedselect3429USEDMULTIPLEselect; end end
  reg [127:0] SR_91;
  wire [127:0] unnamedselect3431USEDMULTIPLEselect;assign unnamedselect3431USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_76):(SR_91)); 
  reg [127:0] unnamedselect3431_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3431_delay1_validunnamednull0_CECE <= unnamedselect3431USEDMULTIPLEselect; end end
  reg [127:0] SR_92;
  wire [127:0] unnamedselect3433USEDMULTIPLEselect;assign unnamedselect3433USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_77):(SR_92)); 
  reg [127:0] unnamedselect3433_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3433_delay1_validunnamednull0_CECE <= unnamedselect3433USEDMULTIPLEselect; end end
  reg [127:0] SR_93;
  wire [127:0] unnamedselect3435USEDMULTIPLEselect;assign unnamedselect3435USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_78):(SR_93)); 
  reg [127:0] unnamedselect3435_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3435_delay1_validunnamednull0_CECE <= unnamedselect3435USEDMULTIPLEselect; end end
  reg [127:0] SR_94;
  wire [127:0] unnamedselect3437USEDMULTIPLEselect;assign unnamedselect3437USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_79):(SR_94)); 
  reg [127:0] unnamedselect3437_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3437_delay1_validunnamednull0_CECE <= unnamedselect3437USEDMULTIPLEselect; end end
  reg [127:0] SR_95;
  wire [127:0] unnamedselect3439USEDMULTIPLEselect;assign unnamedselect3439USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_80):(SR_95)); 
  reg [127:0] unnamedselect3439_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3439_delay1_validunnamednull0_CECE <= unnamedselect3439USEDMULTIPLEselect; end end
  reg [127:0] SR_96;
  wire [127:0] unnamedselect3441USEDMULTIPLEselect;assign unnamedselect3441USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_81):(SR_96)); 
  reg [127:0] unnamedselect3441_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3441_delay1_validunnamednull0_CECE <= unnamedselect3441USEDMULTIPLEselect; end end
  reg [127:0] SR_97;
  wire [127:0] unnamedselect3443USEDMULTIPLEselect;assign unnamedselect3443USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_82):(SR_97)); 
  reg [127:0] unnamedselect3443_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3443_delay1_validunnamednull0_CECE <= unnamedselect3443USEDMULTIPLEselect; end end
  reg [127:0] SR_98;
  wire [127:0] unnamedselect3445USEDMULTIPLEselect;assign unnamedselect3445USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_83):(SR_98)); 
  reg [127:0] unnamedselect3445_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3445_delay1_validunnamednull0_CECE <= unnamedselect3445USEDMULTIPLEselect; end end
  reg [127:0] SR_99;
  wire [127:0] unnamedselect3447USEDMULTIPLEselect;assign unnamedselect3447USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_84):(SR_99)); 
  reg [127:0] unnamedselect3447_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3447_delay1_validunnamednull0_CECE <= unnamedselect3447USEDMULTIPLEselect; end end
  reg [127:0] SR_100;
  wire [127:0] unnamedselect3449USEDMULTIPLEselect;assign unnamedselect3449USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_85):(SR_100)); 
  reg [127:0] unnamedselect3449_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3449_delay1_validunnamednull0_CECE <= unnamedselect3449USEDMULTIPLEselect; end end
  reg [127:0] SR_101;
  wire [127:0] unnamedselect3451USEDMULTIPLEselect;assign unnamedselect3451USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_86):(SR_101)); 
  reg [127:0] unnamedselect3451_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3451_delay1_validunnamednull0_CECE <= unnamedselect3451USEDMULTIPLEselect; end end
  reg [127:0] SR_102;
  wire [127:0] unnamedselect3453USEDMULTIPLEselect;assign unnamedselect3453USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_87):(SR_102)); 
  reg [127:0] unnamedselect3453_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3453_delay1_validunnamednull0_CECE <= unnamedselect3453USEDMULTIPLEselect; end end
  reg [127:0] SR_103;
  wire [127:0] unnamedselect3455USEDMULTIPLEselect;assign unnamedselect3455USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_88):(SR_103)); 
  reg [127:0] unnamedselect3455_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3455_delay1_validunnamednull0_CECE <= unnamedselect3455USEDMULTIPLEselect; end end
  reg [127:0] SR_104;
  wire [127:0] unnamedselect3457USEDMULTIPLEselect;assign unnamedselect3457USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_89):(SR_104)); 
  reg [127:0] unnamedselect3457_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3457_delay1_validunnamednull0_CECE <= unnamedselect3457USEDMULTIPLEselect; end end
  reg [127:0] SR_105;
  wire [127:0] unnamedselect3459USEDMULTIPLEselect;assign unnamedselect3459USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_90):(SR_105)); 
  reg [127:0] unnamedselect3459_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3459_delay1_validunnamednull0_CECE <= unnamedselect3459USEDMULTIPLEselect; end end
  reg [127:0] SR_106;
  wire [127:0] unnamedselect3461USEDMULTIPLEselect;assign unnamedselect3461USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_91):(SR_106)); 
  reg [127:0] unnamedselect3461_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3461_delay1_validunnamednull0_CECE <= unnamedselect3461USEDMULTIPLEselect; end end
  reg [127:0] SR_107;
  wire [127:0] unnamedselect3463USEDMULTIPLEselect;assign unnamedselect3463USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_92):(SR_107)); 
  reg [127:0] unnamedselect3463_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3463_delay1_validunnamednull0_CECE <= unnamedselect3463USEDMULTIPLEselect; end end
  reg [127:0] SR_108;
  wire [127:0] unnamedselect3465USEDMULTIPLEselect;assign unnamedselect3465USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_93):(SR_108)); 
  reg [127:0] unnamedselect3465_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3465_delay1_validunnamednull0_CECE <= unnamedselect3465USEDMULTIPLEselect; end end
  reg [127:0] SR_109;
  wire [127:0] unnamedselect3467USEDMULTIPLEselect;assign unnamedselect3467USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_94):(SR_109)); 
  reg [127:0] unnamedselect3467_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3467_delay1_validunnamednull0_CECE <= unnamedselect3467USEDMULTIPLEselect; end end
  reg [127:0] SR_110;
  wire [127:0] unnamedselect3469USEDMULTIPLEselect;assign unnamedselect3469USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_95):(SR_110)); 
  reg [127:0] unnamedselect3469_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3469_delay1_validunnamednull0_CECE <= unnamedselect3469USEDMULTIPLEselect; end end
  reg [127:0] SR_111;
  wire [127:0] unnamedselect3471USEDMULTIPLEselect;assign unnamedselect3471USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_96):(SR_111)); 
  reg [127:0] unnamedselect3471_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3471_delay1_validunnamednull0_CECE <= unnamedselect3471USEDMULTIPLEselect; end end
  reg [127:0] SR_112;
  wire [127:0] unnamedselect3473USEDMULTIPLEselect;assign unnamedselect3473USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_97):(SR_112)); 
  reg [127:0] unnamedselect3473_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3473_delay1_validunnamednull0_CECE <= unnamedselect3473USEDMULTIPLEselect; end end
  reg [127:0] SR_113;
  wire [127:0] unnamedselect3475USEDMULTIPLEselect;assign unnamedselect3475USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_98):(SR_113)); 
  reg [127:0] unnamedselect3475_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3475_delay1_validunnamednull0_CECE <= unnamedselect3475USEDMULTIPLEselect; end end
  reg [127:0] SR_114;
  wire [127:0] unnamedselect3477USEDMULTIPLEselect;assign unnamedselect3477USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_99):(SR_114)); 
  reg [127:0] unnamedselect3477_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3477_delay1_validunnamednull0_CECE <= unnamedselect3477USEDMULTIPLEselect; end end
  reg [127:0] SR_115;
  wire [127:0] unnamedselect3479USEDMULTIPLEselect;assign unnamedselect3479USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_100):(SR_115)); 
  reg [127:0] unnamedselect3479_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3479_delay1_validunnamednull0_CECE <= unnamedselect3479USEDMULTIPLEselect; end end
  reg [127:0] SR_116;
  wire [127:0] unnamedselect3481USEDMULTIPLEselect;assign unnamedselect3481USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_101):(SR_116)); 
  reg [127:0] unnamedselect3481_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3481_delay1_validunnamednull0_CECE <= unnamedselect3481USEDMULTIPLEselect; end end
  reg [127:0] SR_117;
  wire [127:0] unnamedselect3483USEDMULTIPLEselect;assign unnamedselect3483USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_102):(SR_117)); 
  reg [127:0] unnamedselect3483_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3483_delay1_validunnamednull0_CECE <= unnamedselect3483USEDMULTIPLEselect; end end
  reg [127:0] SR_118;
  wire [127:0] unnamedselect3485USEDMULTIPLEselect;assign unnamedselect3485USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_103):(SR_118)); 
  reg [127:0] unnamedselect3485_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3485_delay1_validunnamednull0_CECE <= unnamedselect3485USEDMULTIPLEselect; end end
  reg [127:0] SR_119;
  wire [127:0] unnamedselect3487USEDMULTIPLEselect;assign unnamedselect3487USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_104):(SR_119)); 
  reg [127:0] unnamedselect3487_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3487_delay1_validunnamednull0_CECE <= unnamedselect3487USEDMULTIPLEselect; end end
  reg [127:0] SR_120;
  wire [127:0] unnamedselect3489USEDMULTIPLEselect;assign unnamedselect3489USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_105):(SR_120)); 
  reg [127:0] unnamedselect3489_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3489_delay1_validunnamednull0_CECE <= unnamedselect3489USEDMULTIPLEselect; end end
  reg [127:0] SR_121;
  wire [127:0] unnamedselect3491USEDMULTIPLEselect;assign unnamedselect3491USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_106):(SR_121)); 
  reg [127:0] unnamedselect3491_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3491_delay1_validunnamednull0_CECE <= unnamedselect3491USEDMULTIPLEselect; end end
  reg [127:0] SR_122;
  wire [127:0] unnamedselect3493USEDMULTIPLEselect;assign unnamedselect3493USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_107):(SR_122)); 
  reg [127:0] unnamedselect3493_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3493_delay1_validunnamednull0_CECE <= unnamedselect3493USEDMULTIPLEselect; end end
  reg [127:0] SR_123;
  wire [127:0] unnamedselect3495USEDMULTIPLEselect;assign unnamedselect3495USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_108):(SR_123)); 
  reg [127:0] unnamedselect3495_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3495_delay1_validunnamednull0_CECE <= unnamedselect3495USEDMULTIPLEselect; end end
  reg [127:0] SR_124;
  wire [127:0] unnamedselect3497USEDMULTIPLEselect;assign unnamedselect3497USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_109):(SR_124)); 
  reg [127:0] unnamedselect3497_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3497_delay1_validunnamednull0_CECE <= unnamedselect3497USEDMULTIPLEselect; end end
  reg [127:0] SR_125;
  wire [127:0] unnamedselect3499USEDMULTIPLEselect;assign unnamedselect3499USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_110):(SR_125)); 
  reg [127:0] unnamedselect3499_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3499_delay1_validunnamednull0_CECE <= unnamedselect3499USEDMULTIPLEselect; end end
  reg [127:0] SR_126;
  wire [127:0] unnamedselect3501USEDMULTIPLEselect;assign unnamedselect3501USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_111):(SR_126)); 
  reg [127:0] unnamedselect3501_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3501_delay1_validunnamednull0_CECE <= unnamedselect3501USEDMULTIPLEselect; end end
  reg [127:0] SR_127;
  wire [127:0] unnamedselect3503USEDMULTIPLEselect;assign unnamedselect3503USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_112):(SR_127)); 
  reg [127:0] unnamedselect3503_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3503_delay1_validunnamednull0_CECE <= unnamedselect3503USEDMULTIPLEselect; end end
  reg [127:0] SR_128;
  wire [127:0] unnamedselect3505USEDMULTIPLEselect;assign unnamedselect3505USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_113):(SR_128)); 
  reg [127:0] unnamedselect3505_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3505_delay1_validunnamednull0_CECE <= unnamedselect3505USEDMULTIPLEselect; end end
  reg [127:0] SR_129;
  wire [127:0] unnamedselect3507USEDMULTIPLEselect;assign unnamedselect3507USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_114):(SR_129)); 
  reg [127:0] unnamedselect3507_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3507_delay1_validunnamednull0_CECE <= unnamedselect3507USEDMULTIPLEselect; end end
  reg [127:0] SR_130;
  wire [127:0] unnamedselect3509USEDMULTIPLEselect;assign unnamedselect3509USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_115):(SR_130)); 
  reg [127:0] unnamedselect3509_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3509_delay1_validunnamednull0_CECE <= unnamedselect3509USEDMULTIPLEselect; end end
  reg [127:0] SR_131;
  wire [127:0] unnamedselect3511USEDMULTIPLEselect;assign unnamedselect3511USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_116):(SR_131)); 
  reg [127:0] unnamedselect3511_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3511_delay1_validunnamednull0_CECE <= unnamedselect3511USEDMULTIPLEselect; end end
  reg [127:0] SR_132;
  wire [127:0] unnamedselect3513USEDMULTIPLEselect;assign unnamedselect3513USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_117):(SR_132)); 
  reg [127:0] unnamedselect3513_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3513_delay1_validunnamednull0_CECE <= unnamedselect3513USEDMULTIPLEselect; end end
  reg [127:0] SR_133;
  wire [127:0] unnamedselect3515USEDMULTIPLEselect;assign unnamedselect3515USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_118):(SR_133)); 
  reg [127:0] unnamedselect3515_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3515_delay1_validunnamednull0_CECE <= unnamedselect3515USEDMULTIPLEselect; end end
  reg [127:0] SR_134;
  wire [127:0] unnamedselect3517USEDMULTIPLEselect;assign unnamedselect3517USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_119):(SR_134)); 
  reg [127:0] unnamedselect3517_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3517_delay1_validunnamednull0_CECE <= unnamedselect3517USEDMULTIPLEselect; end end
  reg [127:0] SR_135;
  wire [127:0] unnamedselect3519USEDMULTIPLEselect;assign unnamedselect3519USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_120):(SR_135)); 
  reg [127:0] unnamedselect3519_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3519_delay1_validunnamednull0_CECE <= unnamedselect3519USEDMULTIPLEselect; end end
  reg [127:0] SR_136;
  wire [127:0] unnamedselect3521USEDMULTIPLEselect;assign unnamedselect3521USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_121):(SR_136)); 
  reg [127:0] unnamedselect3521_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3521_delay1_validunnamednull0_CECE <= unnamedselect3521USEDMULTIPLEselect; end end
  reg [127:0] SR_137;
  wire [127:0] unnamedselect3523USEDMULTIPLEselect;assign unnamedselect3523USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_122):(SR_137)); 
  reg [127:0] unnamedselect3523_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3523_delay1_validunnamednull0_CECE <= unnamedselect3523USEDMULTIPLEselect; end end
  reg [127:0] SR_138;
  wire [127:0] unnamedselect3525USEDMULTIPLEselect;assign unnamedselect3525USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_123):(SR_138)); 
  reg [127:0] unnamedselect3525_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3525_delay1_validunnamednull0_CECE <= unnamedselect3525USEDMULTIPLEselect; end end
  reg [127:0] SR_139;
  wire [127:0] unnamedselect3527USEDMULTIPLEselect;assign unnamedselect3527USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_124):(SR_139)); 
  reg [127:0] unnamedselect3527_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3527_delay1_validunnamednull0_CECE <= unnamedselect3527USEDMULTIPLEselect; end end
  reg [127:0] SR_140;
  wire [127:0] unnamedselect3529USEDMULTIPLEselect;assign unnamedselect3529USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_125):(SR_140)); 
  reg [127:0] unnamedselect3529_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3529_delay1_validunnamednull0_CECE <= unnamedselect3529USEDMULTIPLEselect; end end
  reg [127:0] SR_141;
  wire [127:0] unnamedselect3531USEDMULTIPLEselect;assign unnamedselect3531USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_126):(SR_141)); 
  reg [127:0] unnamedselect3531_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3531_delay1_validunnamednull0_CECE <= unnamedselect3531USEDMULTIPLEselect; end end
  reg [127:0] SR_142;
  wire [127:0] unnamedselect3533USEDMULTIPLEselect;assign unnamedselect3533USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_127):(SR_142)); 
  reg [127:0] unnamedselect3533_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3533_delay1_validunnamednull0_CECE <= unnamedselect3533USEDMULTIPLEselect; end end
  reg [127:0] SR_143;
  wire [127:0] unnamedselect3535USEDMULTIPLEselect;assign unnamedselect3535USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_128):(SR_143)); 
  reg [127:0] unnamedselect3535_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3535_delay1_validunnamednull0_CECE <= unnamedselect3535USEDMULTIPLEselect; end end
  reg [127:0] SR_144;
  wire [127:0] unnamedselect3537USEDMULTIPLEselect;assign unnamedselect3537USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_129):(SR_144)); 
  reg [127:0] unnamedselect3537_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3537_delay1_validunnamednull0_CECE <= unnamedselect3537USEDMULTIPLEselect; end end
  reg [127:0] SR_145;
  wire [127:0] unnamedselect3539USEDMULTIPLEselect;assign unnamedselect3539USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_130):(SR_145)); 
  reg [127:0] unnamedselect3539_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3539_delay1_validunnamednull0_CECE <= unnamedselect3539USEDMULTIPLEselect; end end
  reg [127:0] SR_146;
  wire [127:0] unnamedselect3541USEDMULTIPLEselect;assign unnamedselect3541USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_131):(SR_146)); 
  reg [127:0] unnamedselect3541_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3541_delay1_validunnamednull0_CECE <= unnamedselect3541USEDMULTIPLEselect; end end
  reg [127:0] SR_147;
  wire [127:0] unnamedselect3543USEDMULTIPLEselect;assign unnamedselect3543USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_132):(SR_147)); 
  reg [127:0] unnamedselect3543_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3543_delay1_validunnamednull0_CECE <= unnamedselect3543USEDMULTIPLEselect; end end
  reg [127:0] SR_148;
  wire [127:0] unnamedselect3545USEDMULTIPLEselect;assign unnamedselect3545USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_133):(SR_148)); 
  reg [127:0] unnamedselect3545_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3545_delay1_validunnamednull0_CECE <= unnamedselect3545USEDMULTIPLEselect; end end
  reg [127:0] SR_149;
  wire [127:0] unnamedselect3547USEDMULTIPLEselect;assign unnamedselect3547USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_134):(SR_149)); 
  reg [127:0] unnamedselect3547_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3547_delay1_validunnamednull0_CECE <= unnamedselect3547USEDMULTIPLEselect; end end
  reg [127:0] SR_150;
  wire [127:0] unnamedselect3549USEDMULTIPLEselect;assign unnamedselect3549USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_135):(SR_150)); 
  reg [127:0] unnamedselect3549_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3549_delay1_validunnamednull0_CECE <= unnamedselect3549USEDMULTIPLEselect; end end
  reg [127:0] SR_151;
  wire [127:0] unnamedselect3551USEDMULTIPLEselect;assign unnamedselect3551USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_136):(SR_151)); 
  reg [127:0] unnamedselect3551_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3551_delay1_validunnamednull0_CECE <= unnamedselect3551USEDMULTIPLEselect; end end
  reg [127:0] SR_152;
  wire [127:0] unnamedselect3553USEDMULTIPLEselect;assign unnamedselect3553USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_137):(SR_152)); 
  reg [127:0] unnamedselect3553_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3553_delay1_validunnamednull0_CECE <= unnamedselect3553USEDMULTIPLEselect; end end
  reg [127:0] SR_153;
  wire [127:0] unnamedselect3555USEDMULTIPLEselect;assign unnamedselect3555USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_138):(SR_153)); 
  reg [127:0] unnamedselect3555_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3555_delay1_validunnamednull0_CECE <= unnamedselect3555USEDMULTIPLEselect; end end
  reg [127:0] SR_154;
  wire [127:0] unnamedselect3557USEDMULTIPLEselect;assign unnamedselect3557USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_139):(SR_154)); 
  reg [127:0] unnamedselect3557_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3557_delay1_validunnamednull0_CECE <= unnamedselect3557USEDMULTIPLEselect; end end
  reg [127:0] SR_155;
  wire [127:0] unnamedselect3559USEDMULTIPLEselect;assign unnamedselect3559USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_140):(SR_155)); 
  reg [127:0] unnamedselect3559_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3559_delay1_validunnamednull0_CECE <= unnamedselect3559USEDMULTIPLEselect; end end
  reg [127:0] SR_156;
  wire [127:0] unnamedselect3561USEDMULTIPLEselect;assign unnamedselect3561USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_141):(SR_156)); 
  reg [127:0] unnamedselect3561_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3561_delay1_validunnamednull0_CECE <= unnamedselect3561USEDMULTIPLEselect; end end
  reg [127:0] SR_157;
  wire [127:0] unnamedselect3563USEDMULTIPLEselect;assign unnamedselect3563USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_142):(SR_157)); 
  reg [127:0] unnamedselect3563_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3563_delay1_validunnamednull0_CECE <= unnamedselect3563USEDMULTIPLEselect; end end
  reg [127:0] SR_158;
  wire [127:0] unnamedselect3565USEDMULTIPLEselect;assign unnamedselect3565USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_143):(SR_158)); 
  reg [127:0] unnamedselect3565_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3565_delay1_validunnamednull0_CECE <= unnamedselect3565USEDMULTIPLEselect; end end
  reg [127:0] SR_159;
  wire [127:0] unnamedselect3567USEDMULTIPLEselect;assign unnamedselect3567USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_144):(SR_159)); 
  reg [127:0] unnamedselect3567_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3567_delay1_validunnamednull0_CECE <= unnamedselect3567USEDMULTIPLEselect; end end
  reg [127:0] SR_160;
  wire [127:0] unnamedselect3569USEDMULTIPLEselect;assign unnamedselect3569USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_145):(SR_160)); 
  reg [127:0] unnamedselect3569_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3569_delay1_validunnamednull0_CECE <= unnamedselect3569USEDMULTIPLEselect; end end
  reg [127:0] SR_161;
  wire [127:0] unnamedselect3571USEDMULTIPLEselect;assign unnamedselect3571USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_146):(SR_161)); 
  reg [127:0] unnamedselect3571_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3571_delay1_validunnamednull0_CECE <= unnamedselect3571USEDMULTIPLEselect; end end
  reg [127:0] SR_162;
  wire [127:0] unnamedselect3573USEDMULTIPLEselect;assign unnamedselect3573USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_147):(SR_162)); 
  reg [127:0] unnamedselect3573_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3573_delay1_validunnamednull0_CECE <= unnamedselect3573USEDMULTIPLEselect; end end
  reg [127:0] SR_163;
  wire [127:0] unnamedselect3575USEDMULTIPLEselect;assign unnamedselect3575USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_148):(SR_163)); 
  reg [127:0] unnamedselect3575_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3575_delay1_validunnamednull0_CECE <= unnamedselect3575USEDMULTIPLEselect; end end
  reg [127:0] SR_164;
  wire [127:0] unnamedselect3577USEDMULTIPLEselect;assign unnamedselect3577USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_149):(SR_164)); 
  reg [127:0] unnamedselect3577_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3577_delay1_validunnamednull0_CECE <= unnamedselect3577USEDMULTIPLEselect; end end
  reg [127:0] SR_165;
  wire [127:0] unnamedselect3579USEDMULTIPLEselect;assign unnamedselect3579USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_150):(SR_165)); 
  reg [127:0] unnamedselect3579_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3579_delay1_validunnamednull0_CECE <= unnamedselect3579USEDMULTIPLEselect; end end
  reg [127:0] SR_166;
  wire [127:0] unnamedselect3581USEDMULTIPLEselect;assign unnamedselect3581USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_151):(SR_166)); 
  reg [127:0] unnamedselect3581_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3581_delay1_validunnamednull0_CECE <= unnamedselect3581USEDMULTIPLEselect; end end
  reg [127:0] SR_167;
  wire [127:0] unnamedselect3583USEDMULTIPLEselect;assign unnamedselect3583USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_152):(SR_167)); 
  reg [127:0] unnamedselect3583_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3583_delay1_validunnamednull0_CECE <= unnamedselect3583USEDMULTIPLEselect; end end
  reg [127:0] SR_168;
  wire [127:0] unnamedselect3585USEDMULTIPLEselect;assign unnamedselect3585USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_153):(SR_168)); 
  reg [127:0] unnamedselect3585_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3585_delay1_validunnamednull0_CECE <= unnamedselect3585USEDMULTIPLEselect; end end
  reg [127:0] SR_169;
  wire [127:0] unnamedselect3587USEDMULTIPLEselect;assign unnamedselect3587USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_154):(SR_169)); 
  reg [127:0] unnamedselect3587_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3587_delay1_validunnamednull0_CECE <= unnamedselect3587USEDMULTIPLEselect; end end
  reg [127:0] SR_170;
  wire [127:0] unnamedselect3589USEDMULTIPLEselect;assign unnamedselect3589USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_155):(SR_170)); 
  reg [127:0] unnamedselect3589_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3589_delay1_validunnamednull0_CECE <= unnamedselect3589USEDMULTIPLEselect; end end
  reg [127:0] SR_171;
  wire [127:0] unnamedselect3591USEDMULTIPLEselect;assign unnamedselect3591USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_156):(SR_171)); 
  reg [127:0] unnamedselect3591_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3591_delay1_validunnamednull0_CECE <= unnamedselect3591USEDMULTIPLEselect; end end
  reg [127:0] SR_172;
  wire [127:0] unnamedselect3593USEDMULTIPLEselect;assign unnamedselect3593USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_157):(SR_172)); 
  reg [127:0] unnamedselect3593_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3593_delay1_validunnamednull0_CECE <= unnamedselect3593USEDMULTIPLEselect; end end
  reg [127:0] SR_173;
  wire [127:0] unnamedselect3595USEDMULTIPLEselect;assign unnamedselect3595USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_158):(SR_173)); 
  reg [127:0] unnamedselect3595_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3595_delay1_validunnamednull0_CECE <= unnamedselect3595USEDMULTIPLEselect; end end
  reg [127:0] SR_174;
  wire [127:0] unnamedselect3597USEDMULTIPLEselect;assign unnamedselect3597USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_159):(SR_174)); 
  reg [127:0] unnamedselect3597_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3597_delay1_validunnamednull0_CECE <= unnamedselect3597USEDMULTIPLEselect; end end
  reg [127:0] SR_175;
  wire [127:0] unnamedselect3599USEDMULTIPLEselect;assign unnamedselect3599USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_160):(SR_175)); 
  reg [127:0] unnamedselect3599_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3599_delay1_validunnamednull0_CECE <= unnamedselect3599USEDMULTIPLEselect; end end
  reg [127:0] SR_176;
  wire [127:0] unnamedselect3601USEDMULTIPLEselect;assign unnamedselect3601USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_161):(SR_176)); 
  reg [127:0] unnamedselect3601_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3601_delay1_validunnamednull0_CECE <= unnamedselect3601USEDMULTIPLEselect; end end
  reg [127:0] SR_177;
  wire [127:0] unnamedselect3603USEDMULTIPLEselect;assign unnamedselect3603USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_162):(SR_177)); 
  reg [127:0] unnamedselect3603_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3603_delay1_validunnamednull0_CECE <= unnamedselect3603USEDMULTIPLEselect; end end
  reg [127:0] SR_178;
  wire [127:0] unnamedselect3605USEDMULTIPLEselect;assign unnamedselect3605USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_163):(SR_178)); 
  reg [127:0] unnamedselect3605_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3605_delay1_validunnamednull0_CECE <= unnamedselect3605USEDMULTIPLEselect; end end
  reg [127:0] SR_179;
  wire [127:0] unnamedselect3607USEDMULTIPLEselect;assign unnamedselect3607USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_164):(SR_179)); 
  reg [127:0] unnamedselect3607_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3607_delay1_validunnamednull0_CECE <= unnamedselect3607USEDMULTIPLEselect; end end
  reg [127:0] SR_180;
  wire [127:0] unnamedselect3609USEDMULTIPLEselect;assign unnamedselect3609USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_165):(SR_180)); 
  reg [127:0] unnamedselect3609_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3609_delay1_validunnamednull0_CECE <= unnamedselect3609USEDMULTIPLEselect; end end
  reg [127:0] SR_181;
  wire [127:0] unnamedselect3611USEDMULTIPLEselect;assign unnamedselect3611USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_166):(SR_181)); 
  reg [127:0] unnamedselect3611_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3611_delay1_validunnamednull0_CECE <= unnamedselect3611USEDMULTIPLEselect; end end
  reg [127:0] SR_182;
  wire [127:0] unnamedselect3613USEDMULTIPLEselect;assign unnamedselect3613USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_167):(SR_182)); 
  reg [127:0] unnamedselect3613_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3613_delay1_validunnamednull0_CECE <= unnamedselect3613USEDMULTIPLEselect; end end
  reg [127:0] SR_183;
  wire [127:0] unnamedselect3615USEDMULTIPLEselect;assign unnamedselect3615USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_168):(SR_183)); 
  reg [127:0] unnamedselect3615_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3615_delay1_validunnamednull0_CECE <= unnamedselect3615USEDMULTIPLEselect; end end
  reg [127:0] SR_184;
  wire [127:0] unnamedselect3617USEDMULTIPLEselect;assign unnamedselect3617USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_169):(SR_184)); 
  reg [127:0] unnamedselect3617_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3617_delay1_validunnamednull0_CECE <= unnamedselect3617USEDMULTIPLEselect; end end
  reg [127:0] SR_185;
  wire [127:0] unnamedselect3619USEDMULTIPLEselect;assign unnamedselect3619USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_170):(SR_185)); 
  reg [127:0] unnamedselect3619_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3619_delay1_validunnamednull0_CECE <= unnamedselect3619USEDMULTIPLEselect; end end
  reg [127:0] SR_186;
  wire [127:0] unnamedselect3621USEDMULTIPLEselect;assign unnamedselect3621USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_171):(SR_186)); 
  reg [127:0] unnamedselect3621_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3621_delay1_validunnamednull0_CECE <= unnamedselect3621USEDMULTIPLEselect; end end
  reg [127:0] SR_187;
  wire [127:0] unnamedselect3623USEDMULTIPLEselect;assign unnamedselect3623USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_172):(SR_187)); 
  reg [127:0] unnamedselect3623_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3623_delay1_validunnamednull0_CECE <= unnamedselect3623USEDMULTIPLEselect; end end
  reg [127:0] SR_188;
  wire [127:0] unnamedselect3625USEDMULTIPLEselect;assign unnamedselect3625USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_173):(SR_188)); 
  reg [127:0] unnamedselect3625_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3625_delay1_validunnamednull0_CECE <= unnamedselect3625USEDMULTIPLEselect; end end
  reg [127:0] SR_189;
  wire [127:0] unnamedselect3627USEDMULTIPLEselect;assign unnamedselect3627USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_174):(SR_189)); 
  reg [127:0] unnamedselect3627_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3627_delay1_validunnamednull0_CECE <= unnamedselect3627USEDMULTIPLEselect; end end
  reg [127:0] SR_190;
  wire [127:0] unnamedselect3629USEDMULTIPLEselect;assign unnamedselect3629USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_175):(SR_190)); 
  reg [127:0] unnamedselect3629_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3629_delay1_validunnamednull0_CECE <= unnamedselect3629USEDMULTIPLEselect; end end
  reg [127:0] SR_191;
  wire [127:0] unnamedselect3631USEDMULTIPLEselect;assign unnamedselect3631USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_176):(SR_191)); 
  reg [127:0] unnamedselect3631_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3631_delay1_validunnamednull0_CECE <= unnamedselect3631USEDMULTIPLEselect; end end
  reg [127:0] SR_192;
  wire [127:0] unnamedselect3633USEDMULTIPLEselect;assign unnamedselect3633USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_177):(SR_192)); 
  reg [127:0] unnamedselect3633_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3633_delay1_validunnamednull0_CECE <= unnamedselect3633USEDMULTIPLEselect; end end
  reg [127:0] SR_193;
  wire [127:0] unnamedselect3635USEDMULTIPLEselect;assign unnamedselect3635USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_178):(SR_193)); 
  reg [127:0] unnamedselect3635_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3635_delay1_validunnamednull0_CECE <= unnamedselect3635USEDMULTIPLEselect; end end
  wire [127:0] unnamedselect3637USEDMULTIPLEselect;assign unnamedselect3637USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_179):(SR_194)); 
  reg [127:0] unnamedselect3637_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3637_delay1_validunnamednull0_CECE <= unnamedselect3637USEDMULTIPLEselect; end end
  wire [127:0] unnamedselect3639USEDMULTIPLEselect;assign unnamedselect3639USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_180):(SR_195)); 
  reg [127:0] unnamedselect3639_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3639_delay1_validunnamednull0_CECE <= unnamedselect3639USEDMULTIPLEselect; end end
  wire [127:0] unnamedselect3641USEDMULTIPLEselect;assign unnamedselect3641USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_181):(SR_196)); 
  reg [127:0] unnamedselect3641_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3641_delay1_validunnamednull0_CECE <= unnamedselect3641USEDMULTIPLEselect; end end
  wire [127:0] unnamedselect3643USEDMULTIPLEselect;assign unnamedselect3643USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_182):(SR_197)); 
  reg [127:0] unnamedselect3643_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3643_delay1_validunnamednull0_CECE <= unnamedselect3643USEDMULTIPLEselect; end end
  wire [127:0] unnamedselect3645USEDMULTIPLEselect;assign unnamedselect3645USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_183):(SR_198)); 
  reg [127:0] unnamedselect3645_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3645_delay1_validunnamednull0_CECE <= unnamedselect3645USEDMULTIPLEselect; end end
  wire [127:0] unnamedselect3647USEDMULTIPLEselect;assign unnamedselect3647USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_184):(SR_199)); 
  reg [127:0] unnamedselect3647_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3647_delay1_validunnamednull0_CECE <= unnamedselect3647USEDMULTIPLEselect; end end
  wire [127:0] unnamedselect3649USEDMULTIPLEselect;assign unnamedselect3649USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_185):(SR_200)); 
  reg [127:0] unnamedselect3649_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3649_delay1_validunnamednull0_CECE <= unnamedselect3649USEDMULTIPLEselect; end end
  wire [127:0] unnamedselect3651USEDMULTIPLEselect;assign unnamedselect3651USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_186):(SR_201)); 
  reg [127:0] unnamedselect3651_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3651_delay1_validunnamednull0_CECE <= unnamedselect3651USEDMULTIPLEselect; end end
  wire [127:0] unnamedselect3653USEDMULTIPLEselect;assign unnamedselect3653USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_187):(SR_202)); 
  reg [127:0] unnamedselect3653_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3653_delay1_validunnamednull0_CECE <= unnamedselect3653USEDMULTIPLEselect; end end
  wire [127:0] unnamedselect3655USEDMULTIPLEselect;assign unnamedselect3655USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_188):(SR_203)); 
  reg [127:0] unnamedselect3655_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3655_delay1_validunnamednull0_CECE <= unnamedselect3655USEDMULTIPLEselect; end end
  wire [127:0] unnamedselect3657USEDMULTIPLEselect;assign unnamedselect3657USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_189):(SR_204)); 
  reg [127:0] unnamedselect3657_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3657_delay1_validunnamednull0_CECE <= unnamedselect3657USEDMULTIPLEselect; end end
  wire [127:0] unnamedselect3659USEDMULTIPLEselect;assign unnamedselect3659USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_190):(SR_205)); 
  reg [127:0] unnamedselect3659_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3659_delay1_validunnamednull0_CECE <= unnamedselect3659USEDMULTIPLEselect; end end
  wire [127:0] unnamedselect3661USEDMULTIPLEselect;assign unnamedselect3661USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_191):(SR_206)); 
  reg [127:0] unnamedselect3661_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3661_delay1_validunnamednull0_CECE <= unnamedselect3661USEDMULTIPLEselect; end end
  wire [127:0] unnamedselect3663USEDMULTIPLEselect;assign unnamedselect3663USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(SR_192):(SR_1)); 
  reg [127:0] unnamedselect3663_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3663_delay1_validunnamednull0_CECE <= unnamedselect3663USEDMULTIPLEselect; end end
  wire [127:0] unnamedselect3665USEDMULTIPLEselect;assign unnamedselect3665USEDMULTIPLEselect = ((unnamedbinop2428_readingUSEDMULTIPLEbinop)?(process_input):(SR_2)); 
  reg [127:0] unnamedselect3665_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect3665_delay1_validunnamednull0_CECE <= unnamedselect3665USEDMULTIPLEselect; end end
  reg process_valid_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay1_validunnamednull0_CECE <= process_valid; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_1 <= unnamedselect3255USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_2 <= unnamedselect3257USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_3 <= unnamedselect3259USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_4 <= unnamedselect3261USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_5 <= unnamedselect3263USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_6 <= unnamedselect3265USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_7 <= unnamedselect3267USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_8 <= unnamedselect3269USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_9 <= unnamedselect3271USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_10 <= unnamedselect3273USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_11 <= unnamedselect3275USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_12 <= unnamedselect3277USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_13 <= unnamedselect3279USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_14 <= unnamedselect3281USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_15 <= unnamedselect3283USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_16 <= unnamedselect3285USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_17 <= unnamedselect3287USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_18 <= unnamedselect3289USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_19 <= unnamedselect3291USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_20 <= unnamedselect3293USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_21 <= unnamedselect3295USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_22 <= unnamedselect3297USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_23 <= unnamedselect3299USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_24 <= unnamedselect3301USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_25 <= unnamedselect3303USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_26 <= unnamedselect3305USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_27 <= unnamedselect3307USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_28 <= unnamedselect3309USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_29 <= unnamedselect3311USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_30 <= unnamedselect3313USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_31 <= unnamedselect3315USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_32 <= unnamedselect3317USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_33 <= unnamedselect3319USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_34 <= unnamedselect3321USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_35 <= unnamedselect3323USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_36 <= unnamedselect3325USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_37 <= unnamedselect3327USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_38 <= unnamedselect3329USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_39 <= unnamedselect3331USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_40 <= unnamedselect3333USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_41 <= unnamedselect3335USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_42 <= unnamedselect3337USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_43 <= unnamedselect3339USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_44 <= unnamedselect3341USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_45 <= unnamedselect3343USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_46 <= unnamedselect3345USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_47 <= unnamedselect3347USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_48 <= unnamedselect3349USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_49 <= unnamedselect3351USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_50 <= unnamedselect3353USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_51 <= unnamedselect3355USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_52 <= unnamedselect3357USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_53 <= unnamedselect3359USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_54 <= unnamedselect3361USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_55 <= unnamedselect3363USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_56 <= unnamedselect3365USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_57 <= unnamedselect3367USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_58 <= unnamedselect3369USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_59 <= unnamedselect3371USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_60 <= unnamedselect3373USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_61 <= unnamedselect3375USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_62 <= unnamedselect3377USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_63 <= unnamedselect3379USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_64 <= unnamedselect3381USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_65 <= unnamedselect3383USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_66 <= unnamedselect3385USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_67 <= unnamedselect3387USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_68 <= unnamedselect3389USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_69 <= unnamedselect3391USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_70 <= unnamedselect3393USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_71 <= unnamedselect3395USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_72 <= unnamedselect3397USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_73 <= unnamedselect3399USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_74 <= unnamedselect3401USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_75 <= unnamedselect3403USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_76 <= unnamedselect3405USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_77 <= unnamedselect3407USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_78 <= unnamedselect3409USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_79 <= unnamedselect3411USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_80 <= unnamedselect3413USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_81 <= unnamedselect3415USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_82 <= unnamedselect3417USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_83 <= unnamedselect3419USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_84 <= unnamedselect3421USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_85 <= unnamedselect3423USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_86 <= unnamedselect3425USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_87 <= unnamedselect3427USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_88 <= unnamedselect3429USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_89 <= unnamedselect3431USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_90 <= unnamedselect3433USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_91 <= unnamedselect3435USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_92 <= unnamedselect3437USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_93 <= unnamedselect3439USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_94 <= unnamedselect3441USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_95 <= unnamedselect3443USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_96 <= unnamedselect3445USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_97 <= unnamedselect3447USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_98 <= unnamedselect3449USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_99 <= unnamedselect3451USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_100 <= unnamedselect3453USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_101 <= unnamedselect3455USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_102 <= unnamedselect3457USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_103 <= unnamedselect3459USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_104 <= unnamedselect3461USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_105 <= unnamedselect3463USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_106 <= unnamedselect3465USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_107 <= unnamedselect3467USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_108 <= unnamedselect3469USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_109 <= unnamedselect3471USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_110 <= unnamedselect3473USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_111 <= unnamedselect3475USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_112 <= unnamedselect3477USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_113 <= unnamedselect3479USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_114 <= unnamedselect3481USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_115 <= unnamedselect3483USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_116 <= unnamedselect3485USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_117 <= unnamedselect3487USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_118 <= unnamedselect3489USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_119 <= unnamedselect3491USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_120 <= unnamedselect3493USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_121 <= unnamedselect3495USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_122 <= unnamedselect3497USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_123 <= unnamedselect3499USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_124 <= unnamedselect3501USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_125 <= unnamedselect3503USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_126 <= unnamedselect3505USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_127 <= unnamedselect3507USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_128 <= unnamedselect3509USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_129 <= unnamedselect3511USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_130 <= unnamedselect3513USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_131 <= unnamedselect3515USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_132 <= unnamedselect3517USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_133 <= unnamedselect3519USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_134 <= unnamedselect3521USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_135 <= unnamedselect3523USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_136 <= unnamedselect3525USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_137 <= unnamedselect3527USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_138 <= unnamedselect3529USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_139 <= unnamedselect3531USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_140 <= unnamedselect3533USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_141 <= unnamedselect3535USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_142 <= unnamedselect3537USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_143 <= unnamedselect3539USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_144 <= unnamedselect3541USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_145 <= unnamedselect3543USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_146 <= unnamedselect3545USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_147 <= unnamedselect3547USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_148 <= unnamedselect3549USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_149 <= unnamedselect3551USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_150 <= unnamedselect3553USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_151 <= unnamedselect3555USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_152 <= unnamedselect3557USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_153 <= unnamedselect3559USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_154 <= unnamedselect3561USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_155 <= unnamedselect3563USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_156 <= unnamedselect3565USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_157 <= unnamedselect3567USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_158 <= unnamedselect3569USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_159 <= unnamedselect3571USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_160 <= unnamedselect3573USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_161 <= unnamedselect3575USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_162 <= unnamedselect3577USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_163 <= unnamedselect3579USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_164 <= unnamedselect3581USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_165 <= unnamedselect3583USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_166 <= unnamedselect3585USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_167 <= unnamedselect3587USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_168 <= unnamedselect3589USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_169 <= unnamedselect3591USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_170 <= unnamedselect3593USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_171 <= unnamedselect3595USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_172 <= unnamedselect3597USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_173 <= unnamedselect3599USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_174 <= unnamedselect3601USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_175 <= unnamedselect3603USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_176 <= unnamedselect3605USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_177 <= unnamedselect3607USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_178 <= unnamedselect3609USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_179 <= unnamedselect3611USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_180 <= unnamedselect3613USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_181 <= unnamedselect3615USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_182 <= unnamedselect3617USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_183 <= unnamedselect3619USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_184 <= unnamedselect3621USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_185 <= unnamedselect3623USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_186 <= unnamedselect3625USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_187 <= unnamedselect3627USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_188 <= unnamedselect3629USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_189 <= unnamedselect3631USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_190 <= unnamedselect3633USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_191 <= unnamedselect3635USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_192 <= unnamedselect3637USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_193 <= unnamedselect3639USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_194 <= unnamedselect3641USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_195 <= unnamedselect3643USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_196 <= unnamedselect3645USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_197 <= unnamedselect3647USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_198 <= unnamedselect3649USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_199 <= unnamedselect3651USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_200 <= unnamedselect3653USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_201 <= unnamedselect3655USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_202 <= unnamedselect3657USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_203 <= unnamedselect3659USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_204 <= unnamedselect3661USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_205 <= unnamedselect3663USEDMULTIPLEselect; end end
    always @ (posedge CLK) begin if (process_valid && CE) begin SR_206 <= unnamedselect3665USEDMULTIPLEselect; end end
  wire [15:0] phase_SETBY_OUTPUT;
  assign process_output = {process_valid_delay1_validunnamednull0_CECE,{({unnamedselect3665_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3663_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3661_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3659_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3657_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3655_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3653_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3651_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3649_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3647_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3645_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3643_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3641_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3639_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3637_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3635_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3633_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3631_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3629_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3627_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3625_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3623_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3621_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3619_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3617_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3615_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3613_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3611_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3609_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3607_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3605_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3603_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3601_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3599_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3597_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3595_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3593_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3591_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3589_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3587_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3585_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3583_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3581_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3579_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3577_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3575_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3573_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3571_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3569_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3567_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3565_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3563_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3561_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3559_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3557_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3555_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3553_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3551_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3549_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3547_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3545_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3543_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3541_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3539_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3537_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3535_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3533_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3531_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3529_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3527_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3525_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3523_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3521_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3519_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3517_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3515_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3513_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3511_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3509_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3507_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3505_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3503_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3501_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3499_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3497_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3495_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3493_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3491_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3489_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3487_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3485_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3483_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3481_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3479_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3477_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3475_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3473_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3471_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3469_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3467_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3465_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3463_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3461_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3459_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3457_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3455_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3453_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3451_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3449_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3447_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3445_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3443_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3441_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3439_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3437_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3435_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3433_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3431_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3429_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3427_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3425_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3423_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3421_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3419_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3417_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3415_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3413_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3411_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3409_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3407_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3405_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3403_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3401_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3399_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3397_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3395_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3393_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3391_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3389_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3387_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3385_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3383_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3381_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3379_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3377_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3375_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3373_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3371_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3369_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3367_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3365_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3363_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3361_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3359_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3357_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3355_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3353_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3351_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3349_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3347_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3345_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3343_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3341_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3339_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3337_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3335_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3333_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3331_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3329_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3327_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3325_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3323_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3321_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3319_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3317_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3315_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3313_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3311_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3309_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3307_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3305_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3303_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3301_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3299_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3297_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3295_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3293_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3291_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3289_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3287_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3285_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3283_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3281_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3279_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3277_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3275_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3273_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3271_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3269_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3267_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3265_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3263_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3261_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3259_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3257_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3255_delay1_validunnamednull0_CECE[127:120]}),({unnamedselect3665_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3663_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3661_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3659_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3657_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3655_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3653_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3651_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3649_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3647_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3645_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3643_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3641_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3639_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3637_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3635_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3633_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3631_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3629_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3627_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3625_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3623_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3621_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3619_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3617_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3615_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3613_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3611_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3609_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3607_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3605_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3603_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3601_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3599_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3597_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3595_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3593_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3591_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3589_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3587_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3585_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3583_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3581_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3579_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3577_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3575_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3573_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3571_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3569_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3567_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3565_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3563_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3561_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3559_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3557_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3555_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3553_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3551_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3549_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3547_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3545_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3543_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3541_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3539_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3537_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3535_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3533_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3531_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3529_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3527_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3525_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3523_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3521_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3519_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3517_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3515_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3513_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3511_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3509_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3507_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3505_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3503_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3501_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3499_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3497_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3495_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3493_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3491_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3489_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3487_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3485_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3483_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3481_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3479_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3477_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3475_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3473_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3471_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3469_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3467_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3465_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3463_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3461_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3459_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3457_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3455_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3453_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3451_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3449_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3447_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3445_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3443_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3441_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3439_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3437_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3435_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3433_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3431_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3429_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3427_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3425_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3423_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3421_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3419_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3417_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3415_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3413_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3411_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3409_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3407_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3405_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3403_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3401_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3399_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3397_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3395_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3393_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3391_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3389_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3387_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3385_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3383_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3381_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3379_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3377_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3375_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3373_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3371_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3369_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3367_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3365_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3363_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3361_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3359_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3357_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3355_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3353_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3351_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3349_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3347_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3345_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3343_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3341_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3339_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3337_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3335_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3333_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3331_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3329_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3327_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3325_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3323_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3321_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3319_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3317_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3315_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3313_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3311_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3309_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3307_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3305_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3303_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3301_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3299_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3297_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3295_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3293_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3291_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3289_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3287_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3285_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3283_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3281_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3279_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3277_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3275_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3273_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3271_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3269_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3267_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3265_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3263_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3261_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3259_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3257_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3255_delay1_validunnamednull0_CECE[119:112]}),({unnamedselect3665_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3663_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3661_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3659_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3657_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3655_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3653_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3651_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3649_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3647_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3645_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3643_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3641_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3639_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3637_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3635_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3633_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3631_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3629_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3627_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3625_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3623_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3621_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3619_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3617_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3615_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3613_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3611_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3609_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3607_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3605_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3603_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3601_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3599_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3597_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3595_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3593_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3591_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3589_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3587_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3585_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3583_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3581_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3579_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3577_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3575_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3573_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3571_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3569_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3567_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3565_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3563_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3561_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3559_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3557_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3555_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3553_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3551_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3549_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3547_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3545_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3543_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3541_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3539_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3537_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3535_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3533_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3531_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3529_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3527_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3525_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3523_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3521_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3519_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3517_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3515_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3513_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3511_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3509_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3507_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3505_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3503_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3501_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3499_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3497_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3495_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3493_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3491_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3489_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3487_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3485_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3483_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3481_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3479_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3477_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3475_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3473_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3471_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3469_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3467_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3465_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3463_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3461_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3459_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3457_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3455_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3453_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3451_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3449_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3447_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3445_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3443_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3441_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3439_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3437_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3435_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3433_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3431_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3429_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3427_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3425_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3423_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3421_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3419_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3417_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3415_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3413_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3411_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3409_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3407_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3405_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3403_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3401_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3399_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3397_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3395_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3393_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3391_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3389_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3387_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3385_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3383_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3381_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3379_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3377_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3375_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3373_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3371_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3369_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3367_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3365_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3363_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3361_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3359_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3357_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3355_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3353_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3351_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3349_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3347_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3345_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3343_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3341_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3339_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3337_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3335_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3333_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3331_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3329_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3327_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3325_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3323_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3321_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3319_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3317_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3315_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3313_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3311_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3309_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3307_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3305_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3303_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3301_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3299_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3297_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3295_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3293_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3291_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3289_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3287_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3285_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3283_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3281_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3279_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3277_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3275_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3273_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3271_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3269_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3267_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3265_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3263_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3261_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3259_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3257_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3255_delay1_validunnamednull0_CECE[111:104]}),({unnamedselect3665_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3663_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3661_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3659_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3657_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3655_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3653_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3651_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3649_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3647_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3645_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3643_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3641_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3639_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3637_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3635_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3633_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3631_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3629_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3627_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3625_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3623_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3621_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3619_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3617_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3615_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3613_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3611_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3609_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3607_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3605_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3603_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3601_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3599_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3597_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3595_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3593_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3591_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3589_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3587_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3585_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3583_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3581_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3579_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3577_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3575_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3573_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3571_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3569_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3567_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3565_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3563_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3561_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3559_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3557_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3555_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3553_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3551_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3549_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3547_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3545_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3543_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3541_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3539_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3537_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3535_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3533_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3531_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3529_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3527_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3525_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3523_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3521_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3519_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3517_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3515_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3513_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3511_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3509_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3507_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3505_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3503_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3501_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3499_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3497_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3495_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3493_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3491_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3489_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3487_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3485_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3483_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3481_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3479_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3477_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3475_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3473_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3471_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3469_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3467_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3465_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3463_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3461_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3459_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3457_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3455_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3453_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3451_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3449_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3447_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3445_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3443_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3441_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3439_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3437_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3435_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3433_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3431_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3429_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3427_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3425_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3423_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3421_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3419_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3417_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3415_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3413_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3411_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3409_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3407_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3405_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3403_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3401_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3399_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3397_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3395_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3393_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3391_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3389_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3387_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3385_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3383_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3381_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3379_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3377_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3375_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3373_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3371_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3369_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3367_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3365_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3363_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3361_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3359_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3357_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3355_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3353_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3351_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3349_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3347_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3345_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3343_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3341_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3339_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3337_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3335_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3333_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3331_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3329_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3327_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3325_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3323_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3321_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3319_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3317_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3315_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3313_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3311_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3309_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3307_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3305_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3303_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3301_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3299_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3297_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3295_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3293_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3291_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3289_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3287_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3285_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3283_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3281_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3279_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3277_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3275_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3273_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3271_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3269_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3267_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3265_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3263_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3261_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3259_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3257_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3255_delay1_validunnamednull0_CECE[103:96]}),({unnamedselect3665_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3663_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3661_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3659_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3657_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3655_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3653_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3651_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3649_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3647_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3645_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3643_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3641_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3639_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3637_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3635_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3633_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3631_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3629_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3627_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3625_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3623_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3621_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3619_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3617_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3615_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3613_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3611_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3609_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3607_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3605_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3603_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3601_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3599_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3597_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3595_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3593_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3591_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3589_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3587_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3585_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3583_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3581_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3579_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3577_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3575_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3573_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3571_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3569_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3567_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3565_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3563_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3561_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3559_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3557_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3555_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3553_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3551_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3549_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3547_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3545_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3543_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3541_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3539_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3537_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3535_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3533_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3531_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3529_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3527_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3525_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3523_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3521_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3519_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3517_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3515_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3513_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3511_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3509_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3507_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3505_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3503_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3501_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3499_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3497_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3495_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3493_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3491_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3489_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3487_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3485_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3483_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3481_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3479_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3477_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3475_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3473_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3471_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3469_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3467_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3465_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3463_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3461_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3459_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3457_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3455_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3453_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3451_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3449_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3447_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3445_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3443_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3441_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3439_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3437_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3435_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3433_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3431_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3429_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3427_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3425_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3423_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3421_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3419_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3417_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3415_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3413_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3411_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3409_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3407_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3405_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3403_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3401_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3399_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3397_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3395_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3393_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3391_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3389_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3387_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3385_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3383_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3381_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3379_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3377_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3375_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3373_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3371_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3369_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3367_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3365_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3363_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3361_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3359_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3357_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3355_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3353_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3351_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3349_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3347_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3345_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3343_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3341_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3339_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3337_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3335_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3333_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3331_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3329_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3327_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3325_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3323_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3321_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3319_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3317_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3315_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3313_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3311_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3309_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3307_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3305_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3303_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3301_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3299_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3297_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3295_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3293_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3291_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3289_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3287_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3285_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3283_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3281_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3279_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3277_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3275_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3273_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3271_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3269_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3267_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3265_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3263_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3261_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3259_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3257_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3255_delay1_validunnamednull0_CECE[95:88]}),({unnamedselect3665_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3663_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3661_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3659_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3657_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3655_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3653_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3651_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3649_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3647_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3645_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3643_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3641_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3639_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3637_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3635_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3633_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3631_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3629_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3627_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3625_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3623_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3621_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3619_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3617_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3615_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3613_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3611_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3609_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3607_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3605_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3603_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3601_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3599_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3597_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3595_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3593_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3591_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3589_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3587_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3585_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3583_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3581_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3579_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3577_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3575_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3573_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3571_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3569_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3567_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3565_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3563_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3561_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3559_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3557_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3555_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3553_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3551_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3549_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3547_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3545_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3543_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3541_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3539_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3537_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3535_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3533_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3531_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3529_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3527_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3525_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3523_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3521_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3519_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3517_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3515_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3513_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3511_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3509_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3507_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3505_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3503_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3501_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3499_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3497_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3495_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3493_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3491_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3489_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3487_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3485_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3483_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3481_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3479_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3477_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3475_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3473_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3471_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3469_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3467_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3465_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3463_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3461_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3459_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3457_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3455_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3453_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3451_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3449_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3447_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3445_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3443_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3441_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3439_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3437_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3435_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3433_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3431_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3429_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3427_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3425_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3423_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3421_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3419_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3417_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3415_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3413_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3411_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3409_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3407_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3405_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3403_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3401_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3399_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3397_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3395_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3393_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3391_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3389_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3387_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3385_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3383_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3381_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3379_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3377_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3375_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3373_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3371_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3369_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3367_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3365_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3363_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3361_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3359_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3357_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3355_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3353_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3351_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3349_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3347_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3345_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3343_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3341_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3339_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3337_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3335_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3333_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3331_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3329_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3327_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3325_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3323_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3321_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3319_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3317_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3315_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3313_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3311_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3309_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3307_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3305_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3303_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3301_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3299_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3297_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3295_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3293_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3291_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3289_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3287_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3285_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3283_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3281_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3279_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3277_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3275_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3273_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3271_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3269_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3267_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3265_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3263_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3261_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3259_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3257_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3255_delay1_validunnamednull0_CECE[87:80]}),({unnamedselect3665_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3663_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3661_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3659_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3657_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3655_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3653_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3651_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3649_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3647_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3645_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3643_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3641_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3639_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3637_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3635_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3633_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3631_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3629_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3627_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3625_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3623_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3621_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3619_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3617_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3615_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3613_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3611_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3609_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3607_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3605_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3603_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3601_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3599_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3597_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3595_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3593_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3591_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3589_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3587_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3585_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3583_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3581_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3579_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3577_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3575_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3573_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3571_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3569_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3567_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3565_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3563_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3561_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3559_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3557_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3555_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3553_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3551_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3549_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3547_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3545_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3543_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3541_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3539_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3537_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3535_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3533_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3531_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3529_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3527_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3525_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3523_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3521_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3519_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3517_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3515_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3513_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3511_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3509_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3507_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3505_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3503_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3501_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3499_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3497_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3495_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3493_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3491_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3489_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3487_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3485_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3483_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3481_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3479_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3477_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3475_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3473_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3471_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3469_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3467_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3465_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3463_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3461_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3459_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3457_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3455_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3453_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3451_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3449_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3447_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3445_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3443_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3441_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3439_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3437_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3435_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3433_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3431_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3429_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3427_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3425_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3423_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3421_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3419_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3417_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3415_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3413_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3411_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3409_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3407_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3405_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3403_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3401_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3399_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3397_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3395_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3393_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3391_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3389_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3387_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3385_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3383_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3381_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3379_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3377_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3375_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3373_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3371_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3369_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3367_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3365_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3363_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3361_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3359_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3357_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3355_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3353_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3351_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3349_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3347_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3345_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3343_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3341_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3339_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3337_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3335_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3333_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3331_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3329_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3327_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3325_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3323_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3321_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3319_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3317_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3315_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3313_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3311_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3309_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3307_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3305_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3303_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3301_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3299_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3297_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3295_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3293_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3291_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3289_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3287_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3285_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3283_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3281_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3279_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3277_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3275_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3273_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3271_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3269_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3267_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3265_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3263_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3261_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3259_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3257_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3255_delay1_validunnamednull0_CECE[79:72]}),({unnamedselect3665_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3663_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3661_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3659_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3657_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3655_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3653_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3651_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3649_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3647_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3645_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3643_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3641_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3639_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3637_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3635_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3633_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3631_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3629_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3627_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3625_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3623_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3621_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3619_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3617_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3615_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3613_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3611_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3609_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3607_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3605_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3603_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3601_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3599_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3597_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3595_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3593_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3591_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3589_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3587_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3585_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3583_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3581_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3579_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3577_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3575_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3573_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3571_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3569_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3567_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3565_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3563_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3561_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3559_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3557_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3555_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3553_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3551_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3549_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3547_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3545_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3543_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3541_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3539_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3537_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3535_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3533_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3531_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3529_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3527_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3525_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3523_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3521_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3519_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3517_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3515_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3513_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3511_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3509_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3507_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3505_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3503_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3501_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3499_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3497_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3495_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3493_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3491_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3489_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3487_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3485_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3483_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3481_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3479_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3477_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3475_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3473_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3471_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3469_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3467_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3465_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3463_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3461_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3459_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3457_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3455_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3453_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3451_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3449_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3447_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3445_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3443_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3441_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3439_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3437_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3435_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3433_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3431_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3429_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3427_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3425_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3423_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3421_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3419_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3417_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3415_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3413_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3411_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3409_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3407_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3405_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3403_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3401_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3399_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3397_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3395_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3393_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3391_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3389_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3387_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3385_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3383_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3381_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3379_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3377_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3375_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3373_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3371_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3369_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3367_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3365_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3363_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3361_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3359_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3357_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3355_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3353_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3351_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3349_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3347_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3345_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3343_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3341_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3339_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3337_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3335_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3333_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3331_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3329_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3327_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3325_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3323_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3321_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3319_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3317_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3315_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3313_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3311_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3309_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3307_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3305_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3303_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3301_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3299_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3297_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3295_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3293_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3291_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3289_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3287_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3285_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3283_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3281_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3279_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3277_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3275_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3273_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3271_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3269_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3267_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3265_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3263_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3261_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3259_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3257_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3255_delay1_validunnamednull0_CECE[71:64]}),({unnamedselect3665_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3663_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3661_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3659_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3657_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3655_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3653_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3651_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3649_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3647_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3645_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3643_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3641_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3639_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3637_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3635_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3633_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3631_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3629_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3627_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3625_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3623_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3621_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3619_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3617_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3615_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3613_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3611_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3609_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3607_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3605_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3603_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3601_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3599_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3597_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3595_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3593_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3591_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3589_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3587_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3585_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3583_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3581_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3579_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3577_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3575_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3573_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3571_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3569_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3567_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3565_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3563_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3561_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3559_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3557_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3555_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3553_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3551_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3549_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3547_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3545_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3543_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3541_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3539_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3537_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3535_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3533_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3531_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3529_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3527_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3525_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3523_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3521_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3519_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3517_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3515_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3513_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3511_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3509_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3507_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3505_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3503_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3501_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3499_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3497_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3495_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3493_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3491_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3489_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3487_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3485_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3483_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3481_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3479_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3477_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3475_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3473_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3471_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3469_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3467_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3465_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3463_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3461_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3459_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3457_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3455_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3453_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3451_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3449_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3447_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3445_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3443_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3441_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3439_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3437_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3435_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3433_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3431_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3429_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3427_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3425_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3423_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3421_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3419_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3417_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3415_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3413_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3411_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3409_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3407_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3405_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3403_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3401_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3399_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3397_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3395_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3393_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3391_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3389_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3387_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3385_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3383_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3381_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3379_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3377_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3375_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3373_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3371_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3369_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3367_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3365_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3363_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3361_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3359_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3357_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3355_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3353_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3351_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3349_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3347_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3345_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3343_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3341_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3339_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3337_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3335_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3333_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3331_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3329_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3327_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3325_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3323_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3321_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3319_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3317_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3315_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3313_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3311_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3309_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3307_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3305_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3303_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3301_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3299_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3297_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3295_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3293_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3291_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3289_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3287_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3285_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3283_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3281_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3279_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3277_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3275_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3273_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3271_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3269_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3267_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3265_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3263_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3261_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3259_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3257_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3255_delay1_validunnamednull0_CECE[63:56]}),({unnamedselect3665_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3663_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3661_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3659_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3657_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3655_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3653_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3651_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3649_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3647_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3645_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3643_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3641_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3639_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3637_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3635_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3633_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3631_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3629_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3627_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3625_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3623_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3621_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3619_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3617_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3615_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3613_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3611_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3609_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3607_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3605_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3603_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3601_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3599_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3597_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3595_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3593_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3591_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3589_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3587_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3585_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3583_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3581_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3579_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3577_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3575_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3573_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3571_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3569_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3567_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3565_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3563_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3561_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3559_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3557_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3555_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3553_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3551_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3549_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3547_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3545_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3543_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3541_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3539_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3537_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3535_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3533_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3531_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3529_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3527_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3525_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3523_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3521_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3519_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3517_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3515_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3513_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3511_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3509_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3507_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3505_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3503_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3501_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3499_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3497_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3495_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3493_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3491_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3489_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3487_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3485_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3483_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3481_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3479_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3477_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3475_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3473_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3471_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3469_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3467_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3465_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3463_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3461_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3459_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3457_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3455_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3453_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3451_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3449_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3447_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3445_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3443_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3441_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3439_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3437_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3435_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3433_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3431_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3429_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3427_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3425_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3423_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3421_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3419_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3417_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3415_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3413_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3411_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3409_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3407_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3405_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3403_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3401_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3399_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3397_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3395_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3393_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3391_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3389_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3387_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3385_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3383_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3381_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3379_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3377_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3375_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3373_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3371_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3369_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3367_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3365_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3363_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3361_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3359_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3357_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3355_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3353_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3351_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3349_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3347_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3345_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3343_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3341_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3339_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3337_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3335_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3333_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3331_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3329_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3327_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3325_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3323_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3321_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3319_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3317_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3315_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3313_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3311_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3309_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3307_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3305_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3303_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3301_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3299_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3297_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3295_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3293_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3291_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3289_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3287_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3285_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3283_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3281_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3279_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3277_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3275_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3273_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3271_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3269_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3267_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3265_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3263_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3261_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3259_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3257_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3255_delay1_validunnamednull0_CECE[55:48]}),({unnamedselect3665_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3663_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3661_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3659_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3657_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3655_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3653_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3651_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3649_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3647_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3645_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3643_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3641_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3639_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3637_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3635_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3633_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3631_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3629_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3627_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3625_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3623_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3621_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3619_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3617_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3615_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3613_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3611_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3609_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3607_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3605_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3603_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3601_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3599_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3597_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3595_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3593_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3591_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3589_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3587_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3585_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3583_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3581_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3579_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3577_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3575_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3573_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3571_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3569_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3567_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3565_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3563_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3561_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3559_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3557_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3555_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3553_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3551_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3549_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3547_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3545_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3543_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3541_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3539_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3537_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3535_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3533_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3531_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3529_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3527_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3525_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3523_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3521_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3519_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3517_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3515_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3513_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3511_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3509_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3507_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3505_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3503_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3501_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3499_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3497_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3495_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3493_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3491_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3489_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3487_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3485_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3483_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3481_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3479_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3477_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3475_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3473_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3471_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3469_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3467_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3465_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3463_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3461_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3459_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3457_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3455_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3453_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3451_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3449_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3447_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3445_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3443_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3441_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3439_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3437_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3435_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3433_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3431_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3429_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3427_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3425_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3423_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3421_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3419_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3417_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3415_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3413_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3411_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3409_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3407_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3405_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3403_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3401_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3399_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3397_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3395_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3393_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3391_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3389_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3387_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3385_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3383_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3381_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3379_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3377_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3375_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3373_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3371_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3369_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3367_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3365_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3363_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3361_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3359_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3357_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3355_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3353_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3351_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3349_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3347_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3345_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3343_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3341_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3339_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3337_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3335_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3333_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3331_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3329_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3327_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3325_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3323_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3321_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3319_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3317_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3315_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3313_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3311_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3309_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3307_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3305_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3303_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3301_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3299_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3297_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3295_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3293_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3291_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3289_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3287_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3285_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3283_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3281_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3279_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3277_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3275_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3273_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3271_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3269_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3267_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3265_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3263_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3261_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3259_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3257_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3255_delay1_validunnamednull0_CECE[47:40]}),({unnamedselect3665_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3663_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3661_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3659_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3657_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3655_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3653_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3651_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3649_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3647_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3645_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3643_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3641_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3639_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3637_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3635_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3633_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3631_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3629_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3627_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3625_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3623_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3621_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3619_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3617_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3615_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3613_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3611_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3609_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3607_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3605_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3603_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3601_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3599_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3597_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3595_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3593_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3591_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3589_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3587_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3585_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3583_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3581_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3579_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3577_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3575_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3573_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3571_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3569_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3567_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3565_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3563_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3561_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3559_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3557_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3555_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3553_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3551_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3549_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3547_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3545_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3543_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3541_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3539_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3537_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3535_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3533_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3531_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3529_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3527_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3525_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3523_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3521_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3519_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3517_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3515_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3513_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3511_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3509_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3507_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3505_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3503_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3501_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3499_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3497_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3495_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3493_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3491_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3489_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3487_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3485_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3483_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3481_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3479_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3477_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3475_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3473_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3471_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3469_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3467_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3465_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3463_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3461_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3459_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3457_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3455_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3453_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3451_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3449_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3447_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3445_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3443_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3441_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3439_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3437_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3435_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3433_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3431_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3429_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3427_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3425_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3423_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3421_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3419_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3417_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3415_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3413_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3411_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3409_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3407_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3405_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3403_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3401_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3399_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3397_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3395_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3393_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3391_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3389_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3387_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3385_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3383_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3381_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3379_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3377_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3375_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3373_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3371_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3369_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3367_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3365_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3363_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3361_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3359_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3357_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3355_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3353_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3351_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3349_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3347_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3345_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3343_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3341_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3339_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3337_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3335_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3333_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3331_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3329_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3327_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3325_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3323_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3321_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3319_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3317_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3315_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3313_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3311_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3309_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3307_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3305_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3303_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3301_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3299_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3297_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3295_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3293_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3291_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3289_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3287_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3285_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3283_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3281_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3279_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3277_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3275_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3273_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3271_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3269_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3267_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3265_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3263_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3261_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3259_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3257_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3255_delay1_validunnamednull0_CECE[39:32]}),({unnamedselect3665_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3663_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3661_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3659_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3657_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3655_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3653_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3651_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3649_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3647_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3645_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3643_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3641_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3639_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3637_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3635_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3633_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3631_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3629_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3627_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3625_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3623_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3621_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3619_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3617_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3615_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3613_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3611_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3609_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3607_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3605_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3603_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3601_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3599_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3597_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3595_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3593_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3591_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3589_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3587_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3585_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3583_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3581_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3579_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3577_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3575_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3573_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3571_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3569_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3567_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3565_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3563_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3561_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3559_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3557_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3555_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3553_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3551_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3549_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3547_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3545_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3543_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3541_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3539_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3537_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3535_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3533_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3531_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3529_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3527_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3525_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3523_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3521_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3519_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3517_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3515_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3513_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3511_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3509_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3507_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3505_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3503_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3501_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3499_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3497_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3495_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3493_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3491_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3489_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3487_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3485_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3483_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3481_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3479_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3477_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3475_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3473_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3471_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3469_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3467_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3465_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3463_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3461_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3459_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3457_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3455_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3453_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3451_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3449_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3447_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3445_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3443_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3441_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3439_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3437_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3435_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3433_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3431_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3429_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3427_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3425_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3423_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3421_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3419_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3417_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3415_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3413_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3411_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3409_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3407_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3405_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3403_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3401_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3399_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3397_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3395_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3393_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3391_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3389_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3387_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3385_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3383_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3381_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3379_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3377_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3375_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3373_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3371_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3369_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3367_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3365_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3363_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3361_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3359_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3357_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3355_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3353_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3351_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3349_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3347_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3345_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3343_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3341_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3339_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3337_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3335_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3333_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3331_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3329_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3327_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3325_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3323_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3321_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3319_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3317_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3315_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3313_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3311_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3309_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3307_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3305_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3303_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3301_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3299_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3297_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3295_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3293_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3291_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3289_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3287_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3285_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3283_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3281_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3279_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3277_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3275_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3273_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3271_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3269_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3267_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3265_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3263_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3261_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3259_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3257_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3255_delay1_validunnamednull0_CECE[31:24]}),({unnamedselect3665_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3663_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3661_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3659_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3657_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3655_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3653_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3651_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3649_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3647_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3645_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3643_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3641_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3639_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3637_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3635_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3633_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3631_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3629_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3627_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3625_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3623_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3621_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3619_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3617_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3615_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3613_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3611_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3609_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3607_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3605_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3603_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3601_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3599_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3597_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3595_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3593_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3591_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3589_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3587_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3585_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3583_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3581_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3579_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3577_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3575_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3573_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3571_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3569_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3567_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3565_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3563_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3561_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3559_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3557_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3555_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3553_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3551_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3549_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3547_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3545_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3543_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3541_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3539_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3537_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3535_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3533_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3531_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3529_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3527_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3525_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3523_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3521_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3519_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3517_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3515_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3513_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3511_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3509_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3507_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3505_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3503_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3501_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3499_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3497_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3495_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3493_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3491_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3489_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3487_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3485_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3483_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3481_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3479_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3477_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3475_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3473_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3471_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3469_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3467_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3465_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3463_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3461_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3459_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3457_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3455_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3453_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3451_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3449_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3447_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3445_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3443_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3441_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3439_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3437_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3435_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3433_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3431_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3429_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3427_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3425_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3423_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3421_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3419_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3417_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3415_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3413_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3411_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3409_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3407_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3405_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3403_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3401_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3399_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3397_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3395_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3393_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3391_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3389_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3387_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3385_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3383_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3381_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3379_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3377_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3375_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3373_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3371_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3369_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3367_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3365_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3363_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3361_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3359_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3357_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3355_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3353_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3351_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3349_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3347_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3345_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3343_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3341_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3339_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3337_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3335_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3333_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3331_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3329_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3327_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3325_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3323_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3321_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3319_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3317_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3315_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3313_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3311_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3309_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3307_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3305_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3303_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3301_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3299_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3297_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3295_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3293_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3291_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3289_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3287_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3285_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3283_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3281_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3279_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3277_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3275_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3273_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3271_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3269_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3267_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3265_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3263_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3261_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3259_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3257_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3255_delay1_validunnamednull0_CECE[23:16]}),({unnamedselect3665_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3663_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3661_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3659_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3657_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3655_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3653_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3651_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3649_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3647_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3645_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3643_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3641_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3639_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3637_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3635_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3633_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3631_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3629_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3627_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3625_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3623_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3621_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3619_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3617_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3615_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3613_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3611_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3609_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3607_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3605_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3603_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3601_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3599_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3597_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3595_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3593_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3591_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3589_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3587_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3585_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3583_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3581_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3579_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3577_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3575_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3573_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3571_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3569_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3567_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3565_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3563_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3561_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3559_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3557_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3555_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3553_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3551_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3549_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3547_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3545_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3543_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3541_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3539_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3537_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3535_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3533_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3531_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3529_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3527_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3525_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3523_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3521_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3519_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3517_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3515_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3513_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3511_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3509_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3507_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3505_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3503_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3501_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3499_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3497_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3495_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3493_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3491_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3489_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3487_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3485_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3483_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3481_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3479_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3477_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3475_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3473_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3471_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3469_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3467_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3465_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3463_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3461_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3459_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3457_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3455_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3453_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3451_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3449_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3447_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3445_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3443_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3441_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3439_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3437_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3435_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3433_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3431_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3429_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3427_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3425_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3423_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3421_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3419_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3417_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3415_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3413_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3411_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3409_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3407_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3405_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3403_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3401_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3399_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3397_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3395_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3393_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3391_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3389_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3387_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3385_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3383_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3381_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3379_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3377_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3375_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3373_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3371_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3369_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3367_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3365_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3363_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3361_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3359_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3357_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3355_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3353_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3351_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3349_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3347_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3345_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3343_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3341_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3339_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3337_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3335_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3333_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3331_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3329_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3327_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3325_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3323_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3321_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3319_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3317_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3315_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3313_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3311_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3309_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3307_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3305_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3303_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3301_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3299_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3297_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3295_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3293_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3291_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3289_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3287_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3285_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3283_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3281_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3279_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3277_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3275_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3273_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3271_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3269_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3267_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3265_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3263_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3261_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3259_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3257_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3255_delay1_validunnamednull0_CECE[15:8]}),({unnamedselect3665_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3663_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3661_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3659_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3657_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3655_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3653_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3651_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3649_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3647_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3645_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3643_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3641_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3639_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3637_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3635_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3633_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3631_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3629_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3627_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3625_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3623_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3621_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3619_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3617_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3615_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3613_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3611_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3609_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3607_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3605_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3603_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3601_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3599_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3597_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3595_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3593_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3591_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3589_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3587_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3585_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3583_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3581_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3579_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3577_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3575_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3573_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3571_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3569_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3567_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3565_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3563_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3561_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3559_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3557_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3555_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3553_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3551_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3549_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3547_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3545_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3543_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3541_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3539_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3537_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3535_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3533_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3531_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3529_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3527_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3525_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3523_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3521_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3519_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3517_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3515_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3513_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3511_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3509_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3507_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3505_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3503_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3501_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3499_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3497_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3495_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3493_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3491_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3489_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3487_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3485_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3483_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3481_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3479_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3477_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3475_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3473_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3471_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3469_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3467_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3465_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3463_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3461_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3459_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3457_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3455_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3453_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3451_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3449_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3447_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3445_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3443_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3441_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3439_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3437_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3435_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3433_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3431_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3429_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3427_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3425_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3423_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3421_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3419_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3417_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3415_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3413_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3411_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3409_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3407_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3405_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3403_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3401_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3399_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3397_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3395_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3393_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3391_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3389_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3387_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3385_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3383_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3381_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3379_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3377_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3375_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3373_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3371_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3369_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3367_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3365_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3363_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3361_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3359_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3357_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3355_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3353_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3351_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3349_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3347_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3345_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3343_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3341_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3339_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3337_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3335_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3333_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3331_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3329_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3327_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3325_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3323_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3321_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3319_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3317_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3315_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3313_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3311_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3309_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3307_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3305_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3303_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3301_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3299_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3297_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3295_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3293_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3291_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3289_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3287_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3285_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3283_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3281_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3279_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3277_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3275_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3273_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3271_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3269_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3267_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3265_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3263_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3261_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3259_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3257_delay1_validunnamednull0_CECE[7:0]}),({unnamedselect3255_delay1_validunnamednull0_CECE[7:0]})}};
  // function: ready pure=true delay=0
  // function: reset pure=false delay=0
  // function: process pure=false delay=1
  RegBy_sumwrap_uint16_to7_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_phase"})) phase(.CLK(CLK), .set_valid(reset), .CE(CE), .set_inp((16'd0)), .setby_valid(process_valid), .setby_inp((16'd1)), .SETBY_OUTPUT(phase_SETBY_OUTPUT), .GET_OUTPUT(phase_GET_OUTPUT));
endmodule

module WaitOnInput_SSRPartial_uint8_T0_125(input CLK, output ready, input reset, input CE, input process_valid, input [128:0] process_input, output [26368:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  wire WaitOnInput_inner_ready;
  assign ready = WaitOnInput_inner_ready;
  wire unnamedbinop17307USEDMULTIPLEbinop;assign unnamedbinop17307USEDMULTIPLEbinop = {({({(~WaitOnInput_inner_ready)}||(process_input[128]))}&&process_valid)}; 
  wire [26368:0] WaitOnInput_inner_process_output;
  reg unnamedbinop17307_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedbinop17307_delay1_validunnamednull0_CECE <= unnamedbinop17307USEDMULTIPLEbinop; end end
  assign process_output = {{((WaitOnInput_inner_process_output[26368])&&unnamedbinop17307_delay1_validunnamednull0_CECE)},(WaitOnInput_inner_process_output[26367:0])};
  // function: ready pure=true delay=0
  // function: reset pure=false delay=0
  // function: process pure=false delay=1
  SSRPartial_uint8_T0_125 #(.INSTANCE_NAME({INSTANCE_NAME,"_WaitOnInput_inner"})) WaitOnInput_inner(.CLK(CLK), .ready(WaitOnInput_inner_ready), .reset(reset), .CE(CE), .process_valid(unnamedbinop17307USEDMULTIPLEbinop), .process_input((process_input[127:0])), .process_output(WaitOnInput_inner_process_output));
endmodule

module LiftHandshake_WaitOnInput_SSRPartial_uint8_T0_125(input CLK, input ready_downstream, output ready, input reset, input [128:0] process_input, output [26368:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire inner_WaitOnInput_SSRPartial_uint8_T0_125_ready;
  assign ready = {(inner_WaitOnInput_SSRPartial_uint8_T0_125_ready&&ready_downstream)};
  wire unnamedbinop17341USEDMULTIPLEbinop;assign unnamedbinop17341USEDMULTIPLEbinop = {(reset||ready_downstream)}; 
  wire unnamedunary17342USEDMULTIPLEunary;assign unnamedunary17342USEDMULTIPLEunary = {(~reset)}; 
  wire [26368:0] inner_WaitOnInput_SSRPartial_uint8_T0_125_process_output;
  wire validBitDelay_WaitOnInput_SSRPartial_uint8_T0_125_pushPop_out;
  wire [26368:0] unnamedtuple17352USEDMULTIPLEtuple;assign unnamedtuple17352USEDMULTIPLEtuple = {{((inner_WaitOnInput_SSRPartial_uint8_T0_125_process_output[26368])&&validBitDelay_WaitOnInput_SSRPartial_uint8_T0_125_pushPop_out)},(inner_WaitOnInput_SSRPartial_uint8_T0_125_process_output[26367:0])}; 
  always @(posedge CLK) begin if({(~{((unnamedtuple17352USEDMULTIPLEtuple[26368])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: output valid bit should not be X!",INSTANCE_NAME); end end
  always @(posedge CLK) begin if({(~{((process_input[128])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = unnamedtuple17352USEDMULTIPLEtuple;
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  WaitOnInput_SSRPartial_uint8_T0_125 #(.INSTANCE_NAME({INSTANCE_NAME,"_inner_WaitOnInput_SSRPartial_uint8_T0_125"})) inner_WaitOnInput_SSRPartial_uint8_T0_125(.CLK(CLK), .ready(inner_WaitOnInput_SSRPartial_uint8_T0_125_ready), .reset(reset), .CE(unnamedbinop17341USEDMULTIPLEbinop), .process_valid(unnamedunary17342USEDMULTIPLEunary), .process_input(process_input), .process_output(inner_WaitOnInput_SSRPartial_uint8_T0_125_process_output));
  ShiftRegister_1_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_validBitDelay_WaitOnInput_SSRPartial_uint8_T0_125"})) validBitDelay_WaitOnInput_SSRPartial_uint8_T0_125(.CLK(CLK), .pushPop_valid(unnamedunary17342USEDMULTIPLEunary), .CE(unnamedbinop17341USEDMULTIPLEbinop), .sr_input((1'd1)), .pushPop_out(validBitDelay_WaitOnInput_SSRPartial_uint8_T0_125_pushPop_out), .reset(reset));
endmodule

module slice_typeuint8_206_16__xl0_xh16_yl0_yh15(input CLK, input process_CE, input [26367:0] inp, output [2175:0] process_output);
parameter INSTANCE_NAME="INST";
  assign process_output = {({inp[24855:24848]}),({inp[24847:24840]}),({inp[24839:24832]}),({inp[24831:24824]}),({inp[24823:24816]}),({inp[24815:24808]}),({inp[24807:24800]}),({inp[24799:24792]}),({inp[24791:24784]}),({inp[24783:24776]}),({inp[24775:24768]}),({inp[24767:24760]}),({inp[24759:24752]}),({inp[24751:24744]}),({inp[24743:24736]}),({inp[24735:24728]}),({inp[24727:24720]}),({inp[23207:23200]}),({inp[23199:23192]}),({inp[23191:23184]}),({inp[23183:23176]}),({inp[23175:23168]}),({inp[23167:23160]}),({inp[23159:23152]}),({inp[23151:23144]}),({inp[23143:23136]}),({inp[23135:23128]}),({inp[23127:23120]}),({inp[23119:23112]}),({inp[23111:23104]}),({inp[23103:23096]}),({inp[23095:23088]}),({inp[23087:23080]}),({inp[23079:23072]}),({inp[21559:21552]}),({inp[21551:21544]}),({inp[21543:21536]}),({inp[21535:21528]}),({inp[21527:21520]}),({inp[21519:21512]}),({inp[21511:21504]}),({inp[21503:21496]}),({inp[21495:21488]}),({inp[21487:21480]}),({inp[21479:21472]}),({inp[21471:21464]}),({inp[21463:21456]}),({inp[21455:21448]}),({inp[21447:21440]}),({inp[21439:21432]}),({inp[21431:21424]}),({inp[19911:19904]}),({inp[19903:19896]}),({inp[19895:19888]}),({inp[19887:19880]}),({inp[19879:19872]}),({inp[19871:19864]}),({inp[19863:19856]}),({inp[19855:19848]}),({inp[19847:19840]}),({inp[19839:19832]}),({inp[19831:19824]}),({inp[19823:19816]}),({inp[19815:19808]}),({inp[19807:19800]}),({inp[19799:19792]}),({inp[19791:19784]}),({inp[19783:19776]}),({inp[18263:18256]}),({inp[18255:18248]}),({inp[18247:18240]}),({inp[18239:18232]}),({inp[18231:18224]}),({inp[18223:18216]}),({inp[18215:18208]}),({inp[18207:18200]}),({inp[18199:18192]}),({inp[18191:18184]}),({inp[18183:18176]}),({inp[18175:18168]}),({inp[18167:18160]}),({inp[18159:18152]}),({inp[18151:18144]}),({inp[18143:18136]}),({inp[18135:18128]}),({inp[16615:16608]}),({inp[16607:16600]}),({inp[16599:16592]}),({inp[16591:16584]}),({inp[16583:16576]}),({inp[16575:16568]}),({inp[16567:16560]}),({inp[16559:16552]}),({inp[16551:16544]}),({inp[16543:16536]}),({inp[16535:16528]}),({inp[16527:16520]}),({inp[16519:16512]}),({inp[16511:16504]}),({inp[16503:16496]}),({inp[16495:16488]}),({inp[16487:16480]}),({inp[14967:14960]}),({inp[14959:14952]}),({inp[14951:14944]}),({inp[14943:14936]}),({inp[14935:14928]}),({inp[14927:14920]}),({inp[14919:14912]}),({inp[14911:14904]}),({inp[14903:14896]}),({inp[14895:14888]}),({inp[14887:14880]}),({inp[14879:14872]}),({inp[14871:14864]}),({inp[14863:14856]}),({inp[14855:14848]}),({inp[14847:14840]}),({inp[14839:14832]}),({inp[13319:13312]}),({inp[13311:13304]}),({inp[13303:13296]}),({inp[13295:13288]}),({inp[13287:13280]}),({inp[13279:13272]}),({inp[13271:13264]}),({inp[13263:13256]}),({inp[13255:13248]}),({inp[13247:13240]}),({inp[13239:13232]}),({inp[13231:13224]}),({inp[13223:13216]}),({inp[13215:13208]}),({inp[13207:13200]}),({inp[13199:13192]}),({inp[13191:13184]}),({inp[11671:11664]}),({inp[11663:11656]}),({inp[11655:11648]}),({inp[11647:11640]}),({inp[11639:11632]}),({inp[11631:11624]}),({inp[11623:11616]}),({inp[11615:11608]}),({inp[11607:11600]}),({inp[11599:11592]}),({inp[11591:11584]}),({inp[11583:11576]}),({inp[11575:11568]}),({inp[11567:11560]}),({inp[11559:11552]}),({inp[11551:11544]}),({inp[11543:11536]}),({inp[10023:10016]}),({inp[10015:10008]}),({inp[10007:10000]}),({inp[9999:9992]}),({inp[9991:9984]}),({inp[9983:9976]}),({inp[9975:9968]}),({inp[9967:9960]}),({inp[9959:9952]}),({inp[9951:9944]}),({inp[9943:9936]}),({inp[9935:9928]}),({inp[9927:9920]}),({inp[9919:9912]}),({inp[9911:9904]}),({inp[9903:9896]}),({inp[9895:9888]}),({inp[8375:8368]}),({inp[8367:8360]}),({inp[8359:8352]}),({inp[8351:8344]}),({inp[8343:8336]}),({inp[8335:8328]}),({inp[8327:8320]}),({inp[8319:8312]}),({inp[8311:8304]}),({inp[8303:8296]}),({inp[8295:8288]}),({inp[8287:8280]}),({inp[8279:8272]}),({inp[8271:8264]}),({inp[8263:8256]}),({inp[8255:8248]}),({inp[8247:8240]}),({inp[6727:6720]}),({inp[6719:6712]}),({inp[6711:6704]}),({inp[6703:6696]}),({inp[6695:6688]}),({inp[6687:6680]}),({inp[6679:6672]}),({inp[6671:6664]}),({inp[6663:6656]}),({inp[6655:6648]}),({inp[6647:6640]}),({inp[6639:6632]}),({inp[6631:6624]}),({inp[6623:6616]}),({inp[6615:6608]}),({inp[6607:6600]}),({inp[6599:6592]}),({inp[5079:5072]}),({inp[5071:5064]}),({inp[5063:5056]}),({inp[5055:5048]}),({inp[5047:5040]}),({inp[5039:5032]}),({inp[5031:5024]}),({inp[5023:5016]}),({inp[5015:5008]}),({inp[5007:5000]}),({inp[4999:4992]}),({inp[4991:4984]}),({inp[4983:4976]}),({inp[4975:4968]}),({inp[4967:4960]}),({inp[4959:4952]}),({inp[4951:4944]}),({inp[3431:3424]}),({inp[3423:3416]}),({inp[3415:3408]}),({inp[3407:3400]}),({inp[3399:3392]}),({inp[3391:3384]}),({inp[3383:3376]}),({inp[3375:3368]}),({inp[3367:3360]}),({inp[3359:3352]}),({inp[3351:3344]}),({inp[3343:3336]}),({inp[3335:3328]}),({inp[3327:3320]}),({inp[3319:3312]}),({inp[3311:3304]}),({inp[3303:3296]}),({inp[1783:1776]}),({inp[1775:1768]}),({inp[1767:1760]}),({inp[1759:1752]}),({inp[1751:1744]}),({inp[1743:1736]}),({inp[1735:1728]}),({inp[1727:1720]}),({inp[1719:1712]}),({inp[1711:1704]}),({inp[1703:1696]}),({inp[1695:1688]}),({inp[1687:1680]}),({inp[1679:1672]}),({inp[1671:1664]}),({inp[1663:1656]}),({inp[1655:1648]}),({inp[135:128]}),({inp[127:120]}),({inp[119:112]}),({inp[111:104]}),({inp[103:96]}),({inp[95:88]}),({inp[87:80]}),({inp[79:72]}),({inp[71:64]}),({inp[63:56]}),({inp[55:48]}),({inp[47:40]}),({inp[39:32]}),({inp[31:24]}),({inp[23:16]}),({inp[15:8]}),({inp[7:0]})};
  // function: process pure=true delay=0
endmodule

module MakeHandshake_slice_typeuint8_206_16__xl0_xh16_yl0_yh15(input CLK, input ready_downstream, output ready, input reset, input [26368:0] process_input, output [2176:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  assign ready = ready_downstream;
  wire unnamedbinop18741USEDMULTIPLEbinop;assign unnamedbinop18741USEDMULTIPLEbinop = {(ready_downstream||reset)}; 
  wire unnamedcast18749USEDMULTIPLEcast;assign unnamedcast18749USEDMULTIPLEcast = (process_input[26368]); 
  wire [2175:0] inner_process_output;
  wire validBitDelay_slice_typeuint8_206_16__xl0_xh16_yl0_yh15_pushPop_out;
  always @(posedge CLK) begin if({(~{(unnamedcast18749USEDMULTIPLEcast===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: MakeHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = {validBitDelay_slice_typeuint8_206_16__xl0_xh16_yl0_yh15_pushPop_out,inner_process_output};
  // function: ready pure=true ONLY WIRE
  // function: reset pure=true ONLY WIRE
  // function: process pure=false ONLY WIRE
  ShiftRegister_0_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_validBitDelay_slice_typeuint8_206_16__xl0_xh16_yl0_yh15"})) validBitDelay_slice_typeuint8_206_16__xl0_xh16_yl0_yh15(.CLK(CLK), .CE(unnamedbinop18741USEDMULTIPLEbinop), .sr_input(unnamedcast18749USEDMULTIPLEcast), .pushPop_out(validBitDelay_slice_typeuint8_206_16__xl0_xh16_yl0_yh15_pushPop_out));
  slice_typeuint8_206_16__xl0_xh16_yl0_yh15 #(.INSTANCE_NAME({INSTANCE_NAME,"_inner"})) inner(.CLK(CLK), .process_CE(unnamedbinop18741USEDMULTIPLEbinop), .inp((process_input[26367:0])), .process_output(inner_process_output));
endmodule

module stencilLinebufferPartialOverlap(input CLK, input ready_downstream, output ready, input reset, input [8:0] process_input, output [2176:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire slice_ready;
  wire SSR_ready;
  wire LB_ready;
  assign ready = LB_ready;
  wire [128:0] LB_process_output;
  wire [26368:0] SSR_process_output;
  wire [2176:0] slice_process_output;
  assign process_output = slice_process_output;
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  MakeHandshake_linebuffer_w831_h495_T1_ymin_15_Auint8 #(.INSTANCE_NAME({INSTANCE_NAME,"_LB"})) LB(.CLK(CLK), .ready_downstream(SSR_ready), .ready(LB_ready), .reset(reset), .process_input(process_input), .process_output(LB_process_output));
  LiftHandshake_WaitOnInput_SSRPartial_uint8_T0_125 #(.INSTANCE_NAME({INSTANCE_NAME,"_SSR"})) SSR(.CLK(CLK), .ready_downstream(slice_ready), .ready(SSR_ready), .reset(reset), .process_input(LB_process_output), .process_output(SSR_process_output));
  MakeHandshake_slice_typeuint8_206_16__xl0_xh16_yl0_yh15 #(.INSTANCE_NAME({INSTANCE_NAME,"_slice"})) slice(.CLK(CLK), .ready_downstream(ready_downstream), .ready(slice_ready), .reset(reset), .process_input(SSR_process_output), .process_output(slice_process_output));
endmodule

module unpackStencil_uint8_W16_H16_T2(input CLK, input process_CE, input [2175:0] inp, output [4095:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [7:0] unnamedcast18781USEDMULTIPLEcast;assign unnamedcast18781USEDMULTIPLEcast = ({inp[15:8]}); 
  wire [7:0] unnamedcast18783USEDMULTIPLEcast;assign unnamedcast18783USEDMULTIPLEcast = ({inp[23:16]}); 
  wire [7:0] unnamedcast18785USEDMULTIPLEcast;assign unnamedcast18785USEDMULTIPLEcast = ({inp[31:24]}); 
  wire [7:0] unnamedcast18787USEDMULTIPLEcast;assign unnamedcast18787USEDMULTIPLEcast = ({inp[39:32]}); 
  wire [7:0] unnamedcast18789USEDMULTIPLEcast;assign unnamedcast18789USEDMULTIPLEcast = ({inp[47:40]}); 
  wire [7:0] unnamedcast18791USEDMULTIPLEcast;assign unnamedcast18791USEDMULTIPLEcast = ({inp[55:48]}); 
  wire [7:0] unnamedcast18793USEDMULTIPLEcast;assign unnamedcast18793USEDMULTIPLEcast = ({inp[63:56]}); 
  wire [7:0] unnamedcast18795USEDMULTIPLEcast;assign unnamedcast18795USEDMULTIPLEcast = ({inp[71:64]}); 
  wire [7:0] unnamedcast18797USEDMULTIPLEcast;assign unnamedcast18797USEDMULTIPLEcast = ({inp[79:72]}); 
  wire [7:0] unnamedcast18799USEDMULTIPLEcast;assign unnamedcast18799USEDMULTIPLEcast = ({inp[87:80]}); 
  wire [7:0] unnamedcast18801USEDMULTIPLEcast;assign unnamedcast18801USEDMULTIPLEcast = ({inp[95:88]}); 
  wire [7:0] unnamedcast18803USEDMULTIPLEcast;assign unnamedcast18803USEDMULTIPLEcast = ({inp[103:96]}); 
  wire [7:0] unnamedcast18805USEDMULTIPLEcast;assign unnamedcast18805USEDMULTIPLEcast = ({inp[111:104]}); 
  wire [7:0] unnamedcast18807USEDMULTIPLEcast;assign unnamedcast18807USEDMULTIPLEcast = ({inp[119:112]}); 
  wire [7:0] unnamedcast18809USEDMULTIPLEcast;assign unnamedcast18809USEDMULTIPLEcast = ({inp[127:120]}); 
  wire [7:0] unnamedcast18813USEDMULTIPLEcast;assign unnamedcast18813USEDMULTIPLEcast = ({inp[151:144]}); 
  wire [7:0] unnamedcast18815USEDMULTIPLEcast;assign unnamedcast18815USEDMULTIPLEcast = ({inp[159:152]}); 
  wire [7:0] unnamedcast18817USEDMULTIPLEcast;assign unnamedcast18817USEDMULTIPLEcast = ({inp[167:160]}); 
  wire [7:0] unnamedcast18819USEDMULTIPLEcast;assign unnamedcast18819USEDMULTIPLEcast = ({inp[175:168]}); 
  wire [7:0] unnamedcast18821USEDMULTIPLEcast;assign unnamedcast18821USEDMULTIPLEcast = ({inp[183:176]}); 
  wire [7:0] unnamedcast18823USEDMULTIPLEcast;assign unnamedcast18823USEDMULTIPLEcast = ({inp[191:184]}); 
  wire [7:0] unnamedcast18825USEDMULTIPLEcast;assign unnamedcast18825USEDMULTIPLEcast = ({inp[199:192]}); 
  wire [7:0] unnamedcast18827USEDMULTIPLEcast;assign unnamedcast18827USEDMULTIPLEcast = ({inp[207:200]}); 
  wire [7:0] unnamedcast18829USEDMULTIPLEcast;assign unnamedcast18829USEDMULTIPLEcast = ({inp[215:208]}); 
  wire [7:0] unnamedcast18831USEDMULTIPLEcast;assign unnamedcast18831USEDMULTIPLEcast = ({inp[223:216]}); 
  wire [7:0] unnamedcast18833USEDMULTIPLEcast;assign unnamedcast18833USEDMULTIPLEcast = ({inp[231:224]}); 
  wire [7:0] unnamedcast18835USEDMULTIPLEcast;assign unnamedcast18835USEDMULTIPLEcast = ({inp[239:232]}); 
  wire [7:0] unnamedcast18837USEDMULTIPLEcast;assign unnamedcast18837USEDMULTIPLEcast = ({inp[247:240]}); 
  wire [7:0] unnamedcast18839USEDMULTIPLEcast;assign unnamedcast18839USEDMULTIPLEcast = ({inp[255:248]}); 
  wire [7:0] unnamedcast18841USEDMULTIPLEcast;assign unnamedcast18841USEDMULTIPLEcast = ({inp[263:256]}); 
  wire [7:0] unnamedcast18845USEDMULTIPLEcast;assign unnamedcast18845USEDMULTIPLEcast = ({inp[287:280]}); 
  wire [7:0] unnamedcast18847USEDMULTIPLEcast;assign unnamedcast18847USEDMULTIPLEcast = ({inp[295:288]}); 
  wire [7:0] unnamedcast18849USEDMULTIPLEcast;assign unnamedcast18849USEDMULTIPLEcast = ({inp[303:296]}); 
  wire [7:0] unnamedcast18851USEDMULTIPLEcast;assign unnamedcast18851USEDMULTIPLEcast = ({inp[311:304]}); 
  wire [7:0] unnamedcast18853USEDMULTIPLEcast;assign unnamedcast18853USEDMULTIPLEcast = ({inp[319:312]}); 
  wire [7:0] unnamedcast18855USEDMULTIPLEcast;assign unnamedcast18855USEDMULTIPLEcast = ({inp[327:320]}); 
  wire [7:0] unnamedcast18857USEDMULTIPLEcast;assign unnamedcast18857USEDMULTIPLEcast = ({inp[335:328]}); 
  wire [7:0] unnamedcast18859USEDMULTIPLEcast;assign unnamedcast18859USEDMULTIPLEcast = ({inp[343:336]}); 
  wire [7:0] unnamedcast18861USEDMULTIPLEcast;assign unnamedcast18861USEDMULTIPLEcast = ({inp[351:344]}); 
  wire [7:0] unnamedcast18863USEDMULTIPLEcast;assign unnamedcast18863USEDMULTIPLEcast = ({inp[359:352]}); 
  wire [7:0] unnamedcast18865USEDMULTIPLEcast;assign unnamedcast18865USEDMULTIPLEcast = ({inp[367:360]}); 
  wire [7:0] unnamedcast18867USEDMULTIPLEcast;assign unnamedcast18867USEDMULTIPLEcast = ({inp[375:368]}); 
  wire [7:0] unnamedcast18869USEDMULTIPLEcast;assign unnamedcast18869USEDMULTIPLEcast = ({inp[383:376]}); 
  wire [7:0] unnamedcast18871USEDMULTIPLEcast;assign unnamedcast18871USEDMULTIPLEcast = ({inp[391:384]}); 
  wire [7:0] unnamedcast18873USEDMULTIPLEcast;assign unnamedcast18873USEDMULTIPLEcast = ({inp[399:392]}); 
  wire [7:0] unnamedcast18877USEDMULTIPLEcast;assign unnamedcast18877USEDMULTIPLEcast = ({inp[423:416]}); 
  wire [7:0] unnamedcast18879USEDMULTIPLEcast;assign unnamedcast18879USEDMULTIPLEcast = ({inp[431:424]}); 
  wire [7:0] unnamedcast18881USEDMULTIPLEcast;assign unnamedcast18881USEDMULTIPLEcast = ({inp[439:432]}); 
  wire [7:0] unnamedcast18883USEDMULTIPLEcast;assign unnamedcast18883USEDMULTIPLEcast = ({inp[447:440]}); 
  wire [7:0] unnamedcast18885USEDMULTIPLEcast;assign unnamedcast18885USEDMULTIPLEcast = ({inp[455:448]}); 
  wire [7:0] unnamedcast18887USEDMULTIPLEcast;assign unnamedcast18887USEDMULTIPLEcast = ({inp[463:456]}); 
  wire [7:0] unnamedcast18889USEDMULTIPLEcast;assign unnamedcast18889USEDMULTIPLEcast = ({inp[471:464]}); 
  wire [7:0] unnamedcast18891USEDMULTIPLEcast;assign unnamedcast18891USEDMULTIPLEcast = ({inp[479:472]}); 
  wire [7:0] unnamedcast18893USEDMULTIPLEcast;assign unnamedcast18893USEDMULTIPLEcast = ({inp[487:480]}); 
  wire [7:0] unnamedcast18895USEDMULTIPLEcast;assign unnamedcast18895USEDMULTIPLEcast = ({inp[495:488]}); 
  wire [7:0] unnamedcast18897USEDMULTIPLEcast;assign unnamedcast18897USEDMULTIPLEcast = ({inp[503:496]}); 
  wire [7:0] unnamedcast18899USEDMULTIPLEcast;assign unnamedcast18899USEDMULTIPLEcast = ({inp[511:504]}); 
  wire [7:0] unnamedcast18901USEDMULTIPLEcast;assign unnamedcast18901USEDMULTIPLEcast = ({inp[519:512]}); 
  wire [7:0] unnamedcast18903USEDMULTIPLEcast;assign unnamedcast18903USEDMULTIPLEcast = ({inp[527:520]}); 
  wire [7:0] unnamedcast18905USEDMULTIPLEcast;assign unnamedcast18905USEDMULTIPLEcast = ({inp[535:528]}); 
  wire [7:0] unnamedcast18909USEDMULTIPLEcast;assign unnamedcast18909USEDMULTIPLEcast = ({inp[559:552]}); 
  wire [7:0] unnamedcast18911USEDMULTIPLEcast;assign unnamedcast18911USEDMULTIPLEcast = ({inp[567:560]}); 
  wire [7:0] unnamedcast18913USEDMULTIPLEcast;assign unnamedcast18913USEDMULTIPLEcast = ({inp[575:568]}); 
  wire [7:0] unnamedcast18915USEDMULTIPLEcast;assign unnamedcast18915USEDMULTIPLEcast = ({inp[583:576]}); 
  wire [7:0] unnamedcast18917USEDMULTIPLEcast;assign unnamedcast18917USEDMULTIPLEcast = ({inp[591:584]}); 
  wire [7:0] unnamedcast18919USEDMULTIPLEcast;assign unnamedcast18919USEDMULTIPLEcast = ({inp[599:592]}); 
  wire [7:0] unnamedcast18921USEDMULTIPLEcast;assign unnamedcast18921USEDMULTIPLEcast = ({inp[607:600]}); 
  wire [7:0] unnamedcast18923USEDMULTIPLEcast;assign unnamedcast18923USEDMULTIPLEcast = ({inp[615:608]}); 
  wire [7:0] unnamedcast18925USEDMULTIPLEcast;assign unnamedcast18925USEDMULTIPLEcast = ({inp[623:616]}); 
  wire [7:0] unnamedcast18927USEDMULTIPLEcast;assign unnamedcast18927USEDMULTIPLEcast = ({inp[631:624]}); 
  wire [7:0] unnamedcast18929USEDMULTIPLEcast;assign unnamedcast18929USEDMULTIPLEcast = ({inp[639:632]}); 
  wire [7:0] unnamedcast18931USEDMULTIPLEcast;assign unnamedcast18931USEDMULTIPLEcast = ({inp[647:640]}); 
  wire [7:0] unnamedcast18933USEDMULTIPLEcast;assign unnamedcast18933USEDMULTIPLEcast = ({inp[655:648]}); 
  wire [7:0] unnamedcast18935USEDMULTIPLEcast;assign unnamedcast18935USEDMULTIPLEcast = ({inp[663:656]}); 
  wire [7:0] unnamedcast18937USEDMULTIPLEcast;assign unnamedcast18937USEDMULTIPLEcast = ({inp[671:664]}); 
  wire [7:0] unnamedcast18941USEDMULTIPLEcast;assign unnamedcast18941USEDMULTIPLEcast = ({inp[695:688]}); 
  wire [7:0] unnamedcast18943USEDMULTIPLEcast;assign unnamedcast18943USEDMULTIPLEcast = ({inp[703:696]}); 
  wire [7:0] unnamedcast18945USEDMULTIPLEcast;assign unnamedcast18945USEDMULTIPLEcast = ({inp[711:704]}); 
  wire [7:0] unnamedcast18947USEDMULTIPLEcast;assign unnamedcast18947USEDMULTIPLEcast = ({inp[719:712]}); 
  wire [7:0] unnamedcast18949USEDMULTIPLEcast;assign unnamedcast18949USEDMULTIPLEcast = ({inp[727:720]}); 
  wire [7:0] unnamedcast18951USEDMULTIPLEcast;assign unnamedcast18951USEDMULTIPLEcast = ({inp[735:728]}); 
  wire [7:0] unnamedcast18953USEDMULTIPLEcast;assign unnamedcast18953USEDMULTIPLEcast = ({inp[743:736]}); 
  wire [7:0] unnamedcast18955USEDMULTIPLEcast;assign unnamedcast18955USEDMULTIPLEcast = ({inp[751:744]}); 
  wire [7:0] unnamedcast18957USEDMULTIPLEcast;assign unnamedcast18957USEDMULTIPLEcast = ({inp[759:752]}); 
  wire [7:0] unnamedcast18959USEDMULTIPLEcast;assign unnamedcast18959USEDMULTIPLEcast = ({inp[767:760]}); 
  wire [7:0] unnamedcast18961USEDMULTIPLEcast;assign unnamedcast18961USEDMULTIPLEcast = ({inp[775:768]}); 
  wire [7:0] unnamedcast18963USEDMULTIPLEcast;assign unnamedcast18963USEDMULTIPLEcast = ({inp[783:776]}); 
  wire [7:0] unnamedcast18965USEDMULTIPLEcast;assign unnamedcast18965USEDMULTIPLEcast = ({inp[791:784]}); 
  wire [7:0] unnamedcast18967USEDMULTIPLEcast;assign unnamedcast18967USEDMULTIPLEcast = ({inp[799:792]}); 
  wire [7:0] unnamedcast18969USEDMULTIPLEcast;assign unnamedcast18969USEDMULTIPLEcast = ({inp[807:800]}); 
  wire [7:0] unnamedcast18973USEDMULTIPLEcast;assign unnamedcast18973USEDMULTIPLEcast = ({inp[831:824]}); 
  wire [7:0] unnamedcast18975USEDMULTIPLEcast;assign unnamedcast18975USEDMULTIPLEcast = ({inp[839:832]}); 
  wire [7:0] unnamedcast18977USEDMULTIPLEcast;assign unnamedcast18977USEDMULTIPLEcast = ({inp[847:840]}); 
  wire [7:0] unnamedcast18979USEDMULTIPLEcast;assign unnamedcast18979USEDMULTIPLEcast = ({inp[855:848]}); 
  wire [7:0] unnamedcast18981USEDMULTIPLEcast;assign unnamedcast18981USEDMULTIPLEcast = ({inp[863:856]}); 
  wire [7:0] unnamedcast18983USEDMULTIPLEcast;assign unnamedcast18983USEDMULTIPLEcast = ({inp[871:864]}); 
  wire [7:0] unnamedcast18985USEDMULTIPLEcast;assign unnamedcast18985USEDMULTIPLEcast = ({inp[879:872]}); 
  wire [7:0] unnamedcast18987USEDMULTIPLEcast;assign unnamedcast18987USEDMULTIPLEcast = ({inp[887:880]}); 
  wire [7:0] unnamedcast18989USEDMULTIPLEcast;assign unnamedcast18989USEDMULTIPLEcast = ({inp[895:888]}); 
  wire [7:0] unnamedcast18991USEDMULTIPLEcast;assign unnamedcast18991USEDMULTIPLEcast = ({inp[903:896]}); 
  wire [7:0] unnamedcast18993USEDMULTIPLEcast;assign unnamedcast18993USEDMULTIPLEcast = ({inp[911:904]}); 
  wire [7:0] unnamedcast18995USEDMULTIPLEcast;assign unnamedcast18995USEDMULTIPLEcast = ({inp[919:912]}); 
  wire [7:0] unnamedcast18997USEDMULTIPLEcast;assign unnamedcast18997USEDMULTIPLEcast = ({inp[927:920]}); 
  wire [7:0] unnamedcast18999USEDMULTIPLEcast;assign unnamedcast18999USEDMULTIPLEcast = ({inp[935:928]}); 
  wire [7:0] unnamedcast19001USEDMULTIPLEcast;assign unnamedcast19001USEDMULTIPLEcast = ({inp[943:936]}); 
  wire [7:0] unnamedcast19005USEDMULTIPLEcast;assign unnamedcast19005USEDMULTIPLEcast = ({inp[967:960]}); 
  wire [7:0] unnamedcast19007USEDMULTIPLEcast;assign unnamedcast19007USEDMULTIPLEcast = ({inp[975:968]}); 
  wire [7:0] unnamedcast19009USEDMULTIPLEcast;assign unnamedcast19009USEDMULTIPLEcast = ({inp[983:976]}); 
  wire [7:0] unnamedcast19011USEDMULTIPLEcast;assign unnamedcast19011USEDMULTIPLEcast = ({inp[991:984]}); 
  wire [7:0] unnamedcast19013USEDMULTIPLEcast;assign unnamedcast19013USEDMULTIPLEcast = ({inp[999:992]}); 
  wire [7:0] unnamedcast19015USEDMULTIPLEcast;assign unnamedcast19015USEDMULTIPLEcast = ({inp[1007:1000]}); 
  wire [7:0] unnamedcast19017USEDMULTIPLEcast;assign unnamedcast19017USEDMULTIPLEcast = ({inp[1015:1008]}); 
  wire [7:0] unnamedcast19019USEDMULTIPLEcast;assign unnamedcast19019USEDMULTIPLEcast = ({inp[1023:1016]}); 
  wire [7:0] unnamedcast19021USEDMULTIPLEcast;assign unnamedcast19021USEDMULTIPLEcast = ({inp[1031:1024]}); 
  wire [7:0] unnamedcast19023USEDMULTIPLEcast;assign unnamedcast19023USEDMULTIPLEcast = ({inp[1039:1032]}); 
  wire [7:0] unnamedcast19025USEDMULTIPLEcast;assign unnamedcast19025USEDMULTIPLEcast = ({inp[1047:1040]}); 
  wire [7:0] unnamedcast19027USEDMULTIPLEcast;assign unnamedcast19027USEDMULTIPLEcast = ({inp[1055:1048]}); 
  wire [7:0] unnamedcast19029USEDMULTIPLEcast;assign unnamedcast19029USEDMULTIPLEcast = ({inp[1063:1056]}); 
  wire [7:0] unnamedcast19031USEDMULTIPLEcast;assign unnamedcast19031USEDMULTIPLEcast = ({inp[1071:1064]}); 
  wire [7:0] unnamedcast19033USEDMULTIPLEcast;assign unnamedcast19033USEDMULTIPLEcast = ({inp[1079:1072]}); 
  wire [7:0] unnamedcast19037USEDMULTIPLEcast;assign unnamedcast19037USEDMULTIPLEcast = ({inp[1103:1096]}); 
  wire [7:0] unnamedcast19039USEDMULTIPLEcast;assign unnamedcast19039USEDMULTIPLEcast = ({inp[1111:1104]}); 
  wire [7:0] unnamedcast19041USEDMULTIPLEcast;assign unnamedcast19041USEDMULTIPLEcast = ({inp[1119:1112]}); 
  wire [7:0] unnamedcast19043USEDMULTIPLEcast;assign unnamedcast19043USEDMULTIPLEcast = ({inp[1127:1120]}); 
  wire [7:0] unnamedcast19045USEDMULTIPLEcast;assign unnamedcast19045USEDMULTIPLEcast = ({inp[1135:1128]}); 
  wire [7:0] unnamedcast19047USEDMULTIPLEcast;assign unnamedcast19047USEDMULTIPLEcast = ({inp[1143:1136]}); 
  wire [7:0] unnamedcast19049USEDMULTIPLEcast;assign unnamedcast19049USEDMULTIPLEcast = ({inp[1151:1144]}); 
  wire [7:0] unnamedcast19051USEDMULTIPLEcast;assign unnamedcast19051USEDMULTIPLEcast = ({inp[1159:1152]}); 
  wire [7:0] unnamedcast19053USEDMULTIPLEcast;assign unnamedcast19053USEDMULTIPLEcast = ({inp[1167:1160]}); 
  wire [7:0] unnamedcast19055USEDMULTIPLEcast;assign unnamedcast19055USEDMULTIPLEcast = ({inp[1175:1168]}); 
  wire [7:0] unnamedcast19057USEDMULTIPLEcast;assign unnamedcast19057USEDMULTIPLEcast = ({inp[1183:1176]}); 
  wire [7:0] unnamedcast19059USEDMULTIPLEcast;assign unnamedcast19059USEDMULTIPLEcast = ({inp[1191:1184]}); 
  wire [7:0] unnamedcast19061USEDMULTIPLEcast;assign unnamedcast19061USEDMULTIPLEcast = ({inp[1199:1192]}); 
  wire [7:0] unnamedcast19063USEDMULTIPLEcast;assign unnamedcast19063USEDMULTIPLEcast = ({inp[1207:1200]}); 
  wire [7:0] unnamedcast19065USEDMULTIPLEcast;assign unnamedcast19065USEDMULTIPLEcast = ({inp[1215:1208]}); 
  wire [7:0] unnamedcast19069USEDMULTIPLEcast;assign unnamedcast19069USEDMULTIPLEcast = ({inp[1239:1232]}); 
  wire [7:0] unnamedcast19071USEDMULTIPLEcast;assign unnamedcast19071USEDMULTIPLEcast = ({inp[1247:1240]}); 
  wire [7:0] unnamedcast19073USEDMULTIPLEcast;assign unnamedcast19073USEDMULTIPLEcast = ({inp[1255:1248]}); 
  wire [7:0] unnamedcast19075USEDMULTIPLEcast;assign unnamedcast19075USEDMULTIPLEcast = ({inp[1263:1256]}); 
  wire [7:0] unnamedcast19077USEDMULTIPLEcast;assign unnamedcast19077USEDMULTIPLEcast = ({inp[1271:1264]}); 
  wire [7:0] unnamedcast19079USEDMULTIPLEcast;assign unnamedcast19079USEDMULTIPLEcast = ({inp[1279:1272]}); 
  wire [7:0] unnamedcast19081USEDMULTIPLEcast;assign unnamedcast19081USEDMULTIPLEcast = ({inp[1287:1280]}); 
  wire [7:0] unnamedcast19083USEDMULTIPLEcast;assign unnamedcast19083USEDMULTIPLEcast = ({inp[1295:1288]}); 
  wire [7:0] unnamedcast19085USEDMULTIPLEcast;assign unnamedcast19085USEDMULTIPLEcast = ({inp[1303:1296]}); 
  wire [7:0] unnamedcast19087USEDMULTIPLEcast;assign unnamedcast19087USEDMULTIPLEcast = ({inp[1311:1304]}); 
  wire [7:0] unnamedcast19089USEDMULTIPLEcast;assign unnamedcast19089USEDMULTIPLEcast = ({inp[1319:1312]}); 
  wire [7:0] unnamedcast19091USEDMULTIPLEcast;assign unnamedcast19091USEDMULTIPLEcast = ({inp[1327:1320]}); 
  wire [7:0] unnamedcast19093USEDMULTIPLEcast;assign unnamedcast19093USEDMULTIPLEcast = ({inp[1335:1328]}); 
  wire [7:0] unnamedcast19095USEDMULTIPLEcast;assign unnamedcast19095USEDMULTIPLEcast = ({inp[1343:1336]}); 
  wire [7:0] unnamedcast19097USEDMULTIPLEcast;assign unnamedcast19097USEDMULTIPLEcast = ({inp[1351:1344]}); 
  wire [7:0] unnamedcast19101USEDMULTIPLEcast;assign unnamedcast19101USEDMULTIPLEcast = ({inp[1375:1368]}); 
  wire [7:0] unnamedcast19103USEDMULTIPLEcast;assign unnamedcast19103USEDMULTIPLEcast = ({inp[1383:1376]}); 
  wire [7:0] unnamedcast19105USEDMULTIPLEcast;assign unnamedcast19105USEDMULTIPLEcast = ({inp[1391:1384]}); 
  wire [7:0] unnamedcast19107USEDMULTIPLEcast;assign unnamedcast19107USEDMULTIPLEcast = ({inp[1399:1392]}); 
  wire [7:0] unnamedcast19109USEDMULTIPLEcast;assign unnamedcast19109USEDMULTIPLEcast = ({inp[1407:1400]}); 
  wire [7:0] unnamedcast19111USEDMULTIPLEcast;assign unnamedcast19111USEDMULTIPLEcast = ({inp[1415:1408]}); 
  wire [7:0] unnamedcast19113USEDMULTIPLEcast;assign unnamedcast19113USEDMULTIPLEcast = ({inp[1423:1416]}); 
  wire [7:0] unnamedcast19115USEDMULTIPLEcast;assign unnamedcast19115USEDMULTIPLEcast = ({inp[1431:1424]}); 
  wire [7:0] unnamedcast19117USEDMULTIPLEcast;assign unnamedcast19117USEDMULTIPLEcast = ({inp[1439:1432]}); 
  wire [7:0] unnamedcast19119USEDMULTIPLEcast;assign unnamedcast19119USEDMULTIPLEcast = ({inp[1447:1440]}); 
  wire [7:0] unnamedcast19121USEDMULTIPLEcast;assign unnamedcast19121USEDMULTIPLEcast = ({inp[1455:1448]}); 
  wire [7:0] unnamedcast19123USEDMULTIPLEcast;assign unnamedcast19123USEDMULTIPLEcast = ({inp[1463:1456]}); 
  wire [7:0] unnamedcast19125USEDMULTIPLEcast;assign unnamedcast19125USEDMULTIPLEcast = ({inp[1471:1464]}); 
  wire [7:0] unnamedcast19127USEDMULTIPLEcast;assign unnamedcast19127USEDMULTIPLEcast = ({inp[1479:1472]}); 
  wire [7:0] unnamedcast19129USEDMULTIPLEcast;assign unnamedcast19129USEDMULTIPLEcast = ({inp[1487:1480]}); 
  wire [7:0] unnamedcast19133USEDMULTIPLEcast;assign unnamedcast19133USEDMULTIPLEcast = ({inp[1511:1504]}); 
  wire [7:0] unnamedcast19135USEDMULTIPLEcast;assign unnamedcast19135USEDMULTIPLEcast = ({inp[1519:1512]}); 
  wire [7:0] unnamedcast19137USEDMULTIPLEcast;assign unnamedcast19137USEDMULTIPLEcast = ({inp[1527:1520]}); 
  wire [7:0] unnamedcast19139USEDMULTIPLEcast;assign unnamedcast19139USEDMULTIPLEcast = ({inp[1535:1528]}); 
  wire [7:0] unnamedcast19141USEDMULTIPLEcast;assign unnamedcast19141USEDMULTIPLEcast = ({inp[1543:1536]}); 
  wire [7:0] unnamedcast19143USEDMULTIPLEcast;assign unnamedcast19143USEDMULTIPLEcast = ({inp[1551:1544]}); 
  wire [7:0] unnamedcast19145USEDMULTIPLEcast;assign unnamedcast19145USEDMULTIPLEcast = ({inp[1559:1552]}); 
  wire [7:0] unnamedcast19147USEDMULTIPLEcast;assign unnamedcast19147USEDMULTIPLEcast = ({inp[1567:1560]}); 
  wire [7:0] unnamedcast19149USEDMULTIPLEcast;assign unnamedcast19149USEDMULTIPLEcast = ({inp[1575:1568]}); 
  wire [7:0] unnamedcast19151USEDMULTIPLEcast;assign unnamedcast19151USEDMULTIPLEcast = ({inp[1583:1576]}); 
  wire [7:0] unnamedcast19153USEDMULTIPLEcast;assign unnamedcast19153USEDMULTIPLEcast = ({inp[1591:1584]}); 
  wire [7:0] unnamedcast19155USEDMULTIPLEcast;assign unnamedcast19155USEDMULTIPLEcast = ({inp[1599:1592]}); 
  wire [7:0] unnamedcast19157USEDMULTIPLEcast;assign unnamedcast19157USEDMULTIPLEcast = ({inp[1607:1600]}); 
  wire [7:0] unnamedcast19159USEDMULTIPLEcast;assign unnamedcast19159USEDMULTIPLEcast = ({inp[1615:1608]}); 
  wire [7:0] unnamedcast19161USEDMULTIPLEcast;assign unnamedcast19161USEDMULTIPLEcast = ({inp[1623:1616]}); 
  wire [7:0] unnamedcast19165USEDMULTIPLEcast;assign unnamedcast19165USEDMULTIPLEcast = ({inp[1647:1640]}); 
  wire [7:0] unnamedcast19167USEDMULTIPLEcast;assign unnamedcast19167USEDMULTIPLEcast = ({inp[1655:1648]}); 
  wire [7:0] unnamedcast19169USEDMULTIPLEcast;assign unnamedcast19169USEDMULTIPLEcast = ({inp[1663:1656]}); 
  wire [7:0] unnamedcast19171USEDMULTIPLEcast;assign unnamedcast19171USEDMULTIPLEcast = ({inp[1671:1664]}); 
  wire [7:0] unnamedcast19173USEDMULTIPLEcast;assign unnamedcast19173USEDMULTIPLEcast = ({inp[1679:1672]}); 
  wire [7:0] unnamedcast19175USEDMULTIPLEcast;assign unnamedcast19175USEDMULTIPLEcast = ({inp[1687:1680]}); 
  wire [7:0] unnamedcast19177USEDMULTIPLEcast;assign unnamedcast19177USEDMULTIPLEcast = ({inp[1695:1688]}); 
  wire [7:0] unnamedcast19179USEDMULTIPLEcast;assign unnamedcast19179USEDMULTIPLEcast = ({inp[1703:1696]}); 
  wire [7:0] unnamedcast19181USEDMULTIPLEcast;assign unnamedcast19181USEDMULTIPLEcast = ({inp[1711:1704]}); 
  wire [7:0] unnamedcast19183USEDMULTIPLEcast;assign unnamedcast19183USEDMULTIPLEcast = ({inp[1719:1712]}); 
  wire [7:0] unnamedcast19185USEDMULTIPLEcast;assign unnamedcast19185USEDMULTIPLEcast = ({inp[1727:1720]}); 
  wire [7:0] unnamedcast19187USEDMULTIPLEcast;assign unnamedcast19187USEDMULTIPLEcast = ({inp[1735:1728]}); 
  wire [7:0] unnamedcast19189USEDMULTIPLEcast;assign unnamedcast19189USEDMULTIPLEcast = ({inp[1743:1736]}); 
  wire [7:0] unnamedcast19191USEDMULTIPLEcast;assign unnamedcast19191USEDMULTIPLEcast = ({inp[1751:1744]}); 
  wire [7:0] unnamedcast19193USEDMULTIPLEcast;assign unnamedcast19193USEDMULTIPLEcast = ({inp[1759:1752]}); 
  wire [7:0] unnamedcast19197USEDMULTIPLEcast;assign unnamedcast19197USEDMULTIPLEcast = ({inp[1783:1776]}); 
  wire [7:0] unnamedcast19199USEDMULTIPLEcast;assign unnamedcast19199USEDMULTIPLEcast = ({inp[1791:1784]}); 
  wire [7:0] unnamedcast19201USEDMULTIPLEcast;assign unnamedcast19201USEDMULTIPLEcast = ({inp[1799:1792]}); 
  wire [7:0] unnamedcast19203USEDMULTIPLEcast;assign unnamedcast19203USEDMULTIPLEcast = ({inp[1807:1800]}); 
  wire [7:0] unnamedcast19205USEDMULTIPLEcast;assign unnamedcast19205USEDMULTIPLEcast = ({inp[1815:1808]}); 
  wire [7:0] unnamedcast19207USEDMULTIPLEcast;assign unnamedcast19207USEDMULTIPLEcast = ({inp[1823:1816]}); 
  wire [7:0] unnamedcast19209USEDMULTIPLEcast;assign unnamedcast19209USEDMULTIPLEcast = ({inp[1831:1824]}); 
  wire [7:0] unnamedcast19211USEDMULTIPLEcast;assign unnamedcast19211USEDMULTIPLEcast = ({inp[1839:1832]}); 
  wire [7:0] unnamedcast19213USEDMULTIPLEcast;assign unnamedcast19213USEDMULTIPLEcast = ({inp[1847:1840]}); 
  wire [7:0] unnamedcast19215USEDMULTIPLEcast;assign unnamedcast19215USEDMULTIPLEcast = ({inp[1855:1848]}); 
  wire [7:0] unnamedcast19217USEDMULTIPLEcast;assign unnamedcast19217USEDMULTIPLEcast = ({inp[1863:1856]}); 
  wire [7:0] unnamedcast19219USEDMULTIPLEcast;assign unnamedcast19219USEDMULTIPLEcast = ({inp[1871:1864]}); 
  wire [7:0] unnamedcast19221USEDMULTIPLEcast;assign unnamedcast19221USEDMULTIPLEcast = ({inp[1879:1872]}); 
  wire [7:0] unnamedcast19223USEDMULTIPLEcast;assign unnamedcast19223USEDMULTIPLEcast = ({inp[1887:1880]}); 
  wire [7:0] unnamedcast19225USEDMULTIPLEcast;assign unnamedcast19225USEDMULTIPLEcast = ({inp[1895:1888]}); 
  wire [7:0] unnamedcast19229USEDMULTIPLEcast;assign unnamedcast19229USEDMULTIPLEcast = ({inp[1919:1912]}); 
  wire [7:0] unnamedcast19231USEDMULTIPLEcast;assign unnamedcast19231USEDMULTIPLEcast = ({inp[1927:1920]}); 
  wire [7:0] unnamedcast19233USEDMULTIPLEcast;assign unnamedcast19233USEDMULTIPLEcast = ({inp[1935:1928]}); 
  wire [7:0] unnamedcast19235USEDMULTIPLEcast;assign unnamedcast19235USEDMULTIPLEcast = ({inp[1943:1936]}); 
  wire [7:0] unnamedcast19237USEDMULTIPLEcast;assign unnamedcast19237USEDMULTIPLEcast = ({inp[1951:1944]}); 
  wire [7:0] unnamedcast19239USEDMULTIPLEcast;assign unnamedcast19239USEDMULTIPLEcast = ({inp[1959:1952]}); 
  wire [7:0] unnamedcast19241USEDMULTIPLEcast;assign unnamedcast19241USEDMULTIPLEcast = ({inp[1967:1960]}); 
  wire [7:0] unnamedcast19243USEDMULTIPLEcast;assign unnamedcast19243USEDMULTIPLEcast = ({inp[1975:1968]}); 
  wire [7:0] unnamedcast19245USEDMULTIPLEcast;assign unnamedcast19245USEDMULTIPLEcast = ({inp[1983:1976]}); 
  wire [7:0] unnamedcast19247USEDMULTIPLEcast;assign unnamedcast19247USEDMULTIPLEcast = ({inp[1991:1984]}); 
  wire [7:0] unnamedcast19249USEDMULTIPLEcast;assign unnamedcast19249USEDMULTIPLEcast = ({inp[1999:1992]}); 
  wire [7:0] unnamedcast19251USEDMULTIPLEcast;assign unnamedcast19251USEDMULTIPLEcast = ({inp[2007:2000]}); 
  wire [7:0] unnamedcast19253USEDMULTIPLEcast;assign unnamedcast19253USEDMULTIPLEcast = ({inp[2015:2008]}); 
  wire [7:0] unnamedcast19255USEDMULTIPLEcast;assign unnamedcast19255USEDMULTIPLEcast = ({inp[2023:2016]}); 
  wire [7:0] unnamedcast19257USEDMULTIPLEcast;assign unnamedcast19257USEDMULTIPLEcast = ({inp[2031:2024]}); 
  wire [7:0] unnamedcast19261USEDMULTIPLEcast;assign unnamedcast19261USEDMULTIPLEcast = ({inp[2055:2048]}); 
  wire [7:0] unnamedcast19263USEDMULTIPLEcast;assign unnamedcast19263USEDMULTIPLEcast = ({inp[2063:2056]}); 
  wire [7:0] unnamedcast19265USEDMULTIPLEcast;assign unnamedcast19265USEDMULTIPLEcast = ({inp[2071:2064]}); 
  wire [7:0] unnamedcast19267USEDMULTIPLEcast;assign unnamedcast19267USEDMULTIPLEcast = ({inp[2079:2072]}); 
  wire [7:0] unnamedcast19269USEDMULTIPLEcast;assign unnamedcast19269USEDMULTIPLEcast = ({inp[2087:2080]}); 
  wire [7:0] unnamedcast19271USEDMULTIPLEcast;assign unnamedcast19271USEDMULTIPLEcast = ({inp[2095:2088]}); 
  wire [7:0] unnamedcast19273USEDMULTIPLEcast;assign unnamedcast19273USEDMULTIPLEcast = ({inp[2103:2096]}); 
  wire [7:0] unnamedcast19275USEDMULTIPLEcast;assign unnamedcast19275USEDMULTIPLEcast = ({inp[2111:2104]}); 
  wire [7:0] unnamedcast19277USEDMULTIPLEcast;assign unnamedcast19277USEDMULTIPLEcast = ({inp[2119:2112]}); 
  wire [7:0] unnamedcast19279USEDMULTIPLEcast;assign unnamedcast19279USEDMULTIPLEcast = ({inp[2127:2120]}); 
  wire [7:0] unnamedcast19281USEDMULTIPLEcast;assign unnamedcast19281USEDMULTIPLEcast = ({inp[2135:2128]}); 
  wire [7:0] unnamedcast19283USEDMULTIPLEcast;assign unnamedcast19283USEDMULTIPLEcast = ({inp[2143:2136]}); 
  wire [7:0] unnamedcast19285USEDMULTIPLEcast;assign unnamedcast19285USEDMULTIPLEcast = ({inp[2151:2144]}); 
  wire [7:0] unnamedcast19287USEDMULTIPLEcast;assign unnamedcast19287USEDMULTIPLEcast = ({inp[2159:2152]}); 
  wire [7:0] unnamedcast19289USEDMULTIPLEcast;assign unnamedcast19289USEDMULTIPLEcast = ({inp[2167:2160]}); 
  assign process_output = {{({inp[2175:2168]}),unnamedcast19289USEDMULTIPLEcast,unnamedcast19287USEDMULTIPLEcast,unnamedcast19285USEDMULTIPLEcast,unnamedcast19283USEDMULTIPLEcast,unnamedcast19281USEDMULTIPLEcast,unnamedcast19279USEDMULTIPLEcast,unnamedcast19277USEDMULTIPLEcast,unnamedcast19275USEDMULTIPLEcast,unnamedcast19273USEDMULTIPLEcast,unnamedcast19271USEDMULTIPLEcast,unnamedcast19269USEDMULTIPLEcast,unnamedcast19267USEDMULTIPLEcast,unnamedcast19265USEDMULTIPLEcast,unnamedcast19263USEDMULTIPLEcast,unnamedcast19261USEDMULTIPLEcast,({inp[2039:2032]}),unnamedcast19257USEDMULTIPLEcast,unnamedcast19255USEDMULTIPLEcast,unnamedcast19253USEDMULTIPLEcast,unnamedcast19251USEDMULTIPLEcast,unnamedcast19249USEDMULTIPLEcast,unnamedcast19247USEDMULTIPLEcast,unnamedcast19245USEDMULTIPLEcast,unnamedcast19243USEDMULTIPLEcast,unnamedcast19241USEDMULTIPLEcast,unnamedcast19239USEDMULTIPLEcast,unnamedcast19237USEDMULTIPLEcast,unnamedcast19235USEDMULTIPLEcast,unnamedcast19233USEDMULTIPLEcast,unnamedcast19231USEDMULTIPLEcast,unnamedcast19229USEDMULTIPLEcast,({inp[1903:1896]}),unnamedcast19225USEDMULTIPLEcast,unnamedcast19223USEDMULTIPLEcast,unnamedcast19221USEDMULTIPLEcast,unnamedcast19219USEDMULTIPLEcast,unnamedcast19217USEDMULTIPLEcast,unnamedcast19215USEDMULTIPLEcast,unnamedcast19213USEDMULTIPLEcast,unnamedcast19211USEDMULTIPLEcast,unnamedcast19209USEDMULTIPLEcast,unnamedcast19207USEDMULTIPLEcast,unnamedcast19205USEDMULTIPLEcast,unnamedcast19203USEDMULTIPLEcast,unnamedcast19201USEDMULTIPLEcast,unnamedcast19199USEDMULTIPLEcast,unnamedcast19197USEDMULTIPLEcast,({inp[1767:1760]}),unnamedcast19193USEDMULTIPLEcast,unnamedcast19191USEDMULTIPLEcast,unnamedcast19189USEDMULTIPLEcast,unnamedcast19187USEDMULTIPLEcast,unnamedcast19185USEDMULTIPLEcast,unnamedcast19183USEDMULTIPLEcast,unnamedcast19181USEDMULTIPLEcast,unnamedcast19179USEDMULTIPLEcast,unnamedcast19177USEDMULTIPLEcast,unnamedcast19175USEDMULTIPLEcast,unnamedcast19173USEDMULTIPLEcast,unnamedcast19171USEDMULTIPLEcast,unnamedcast19169USEDMULTIPLEcast,unnamedcast19167USEDMULTIPLEcast,unnamedcast19165USEDMULTIPLEcast,({inp[1631:1624]}),unnamedcast19161USEDMULTIPLEcast,unnamedcast19159USEDMULTIPLEcast,unnamedcast19157USEDMULTIPLEcast,unnamedcast19155USEDMULTIPLEcast,unnamedcast19153USEDMULTIPLEcast,unnamedcast19151USEDMULTIPLEcast,unnamedcast19149USEDMULTIPLEcast,unnamedcast19147USEDMULTIPLEcast,unnamedcast19145USEDMULTIPLEcast,unnamedcast19143USEDMULTIPLEcast,unnamedcast19141USEDMULTIPLEcast,unnamedcast19139USEDMULTIPLEcast,unnamedcast19137USEDMULTIPLEcast,unnamedcast19135USEDMULTIPLEcast,unnamedcast19133USEDMULTIPLEcast,({inp[1495:1488]}),unnamedcast19129USEDMULTIPLEcast,unnamedcast19127USEDMULTIPLEcast,unnamedcast19125USEDMULTIPLEcast,unnamedcast19123USEDMULTIPLEcast,unnamedcast19121USEDMULTIPLEcast,unnamedcast19119USEDMULTIPLEcast,unnamedcast19117USEDMULTIPLEcast,unnamedcast19115USEDMULTIPLEcast,unnamedcast19113USEDMULTIPLEcast,unnamedcast19111USEDMULTIPLEcast,unnamedcast19109USEDMULTIPLEcast,unnamedcast19107USEDMULTIPLEcast,unnamedcast19105USEDMULTIPLEcast,unnamedcast19103USEDMULTIPLEcast,unnamedcast19101USEDMULTIPLEcast,({inp[1359:1352]}),unnamedcast19097USEDMULTIPLEcast,unnamedcast19095USEDMULTIPLEcast,unnamedcast19093USEDMULTIPLEcast,unnamedcast19091USEDMULTIPLEcast,unnamedcast19089USEDMULTIPLEcast,unnamedcast19087USEDMULTIPLEcast,unnamedcast19085USEDMULTIPLEcast,unnamedcast19083USEDMULTIPLEcast,unnamedcast19081USEDMULTIPLEcast,unnamedcast19079USEDMULTIPLEcast,unnamedcast19077USEDMULTIPLEcast,unnamedcast19075USEDMULTIPLEcast,unnamedcast19073USEDMULTIPLEcast,unnamedcast19071USEDMULTIPLEcast,unnamedcast19069USEDMULTIPLEcast,({inp[1223:1216]}),unnamedcast19065USEDMULTIPLEcast,unnamedcast19063USEDMULTIPLEcast,unnamedcast19061USEDMULTIPLEcast,unnamedcast19059USEDMULTIPLEcast,unnamedcast19057USEDMULTIPLEcast,unnamedcast19055USEDMULTIPLEcast,unnamedcast19053USEDMULTIPLEcast,unnamedcast19051USEDMULTIPLEcast,unnamedcast19049USEDMULTIPLEcast,unnamedcast19047USEDMULTIPLEcast,unnamedcast19045USEDMULTIPLEcast,unnamedcast19043USEDMULTIPLEcast,unnamedcast19041USEDMULTIPLEcast,unnamedcast19039USEDMULTIPLEcast,unnamedcast19037USEDMULTIPLEcast,({inp[1087:1080]}),unnamedcast19033USEDMULTIPLEcast,unnamedcast19031USEDMULTIPLEcast,unnamedcast19029USEDMULTIPLEcast,unnamedcast19027USEDMULTIPLEcast,unnamedcast19025USEDMULTIPLEcast,unnamedcast19023USEDMULTIPLEcast,unnamedcast19021USEDMULTIPLEcast,unnamedcast19019USEDMULTIPLEcast,unnamedcast19017USEDMULTIPLEcast,unnamedcast19015USEDMULTIPLEcast,unnamedcast19013USEDMULTIPLEcast,unnamedcast19011USEDMULTIPLEcast,unnamedcast19009USEDMULTIPLEcast,unnamedcast19007USEDMULTIPLEcast,unnamedcast19005USEDMULTIPLEcast,({inp[951:944]}),unnamedcast19001USEDMULTIPLEcast,unnamedcast18999USEDMULTIPLEcast,unnamedcast18997USEDMULTIPLEcast,unnamedcast18995USEDMULTIPLEcast,unnamedcast18993USEDMULTIPLEcast,unnamedcast18991USEDMULTIPLEcast,unnamedcast18989USEDMULTIPLEcast,unnamedcast18987USEDMULTIPLEcast,unnamedcast18985USEDMULTIPLEcast,unnamedcast18983USEDMULTIPLEcast,unnamedcast18981USEDMULTIPLEcast,unnamedcast18979USEDMULTIPLEcast,unnamedcast18977USEDMULTIPLEcast,unnamedcast18975USEDMULTIPLEcast,unnamedcast18973USEDMULTIPLEcast,({inp[815:808]}),unnamedcast18969USEDMULTIPLEcast,unnamedcast18967USEDMULTIPLEcast,unnamedcast18965USEDMULTIPLEcast,unnamedcast18963USEDMULTIPLEcast,unnamedcast18961USEDMULTIPLEcast,unnamedcast18959USEDMULTIPLEcast,unnamedcast18957USEDMULTIPLEcast,unnamedcast18955USEDMULTIPLEcast,unnamedcast18953USEDMULTIPLEcast,unnamedcast18951USEDMULTIPLEcast,unnamedcast18949USEDMULTIPLEcast,unnamedcast18947USEDMULTIPLEcast,unnamedcast18945USEDMULTIPLEcast,unnamedcast18943USEDMULTIPLEcast,unnamedcast18941USEDMULTIPLEcast,({inp[679:672]}),unnamedcast18937USEDMULTIPLEcast,unnamedcast18935USEDMULTIPLEcast,unnamedcast18933USEDMULTIPLEcast,unnamedcast18931USEDMULTIPLEcast,unnamedcast18929USEDMULTIPLEcast,unnamedcast18927USEDMULTIPLEcast,unnamedcast18925USEDMULTIPLEcast,unnamedcast18923USEDMULTIPLEcast,unnamedcast18921USEDMULTIPLEcast,unnamedcast18919USEDMULTIPLEcast,unnamedcast18917USEDMULTIPLEcast,unnamedcast18915USEDMULTIPLEcast,unnamedcast18913USEDMULTIPLEcast,unnamedcast18911USEDMULTIPLEcast,unnamedcast18909USEDMULTIPLEcast,({inp[543:536]}),unnamedcast18905USEDMULTIPLEcast,unnamedcast18903USEDMULTIPLEcast,unnamedcast18901USEDMULTIPLEcast,unnamedcast18899USEDMULTIPLEcast,unnamedcast18897USEDMULTIPLEcast,unnamedcast18895USEDMULTIPLEcast,unnamedcast18893USEDMULTIPLEcast,unnamedcast18891USEDMULTIPLEcast,unnamedcast18889USEDMULTIPLEcast,unnamedcast18887USEDMULTIPLEcast,unnamedcast18885USEDMULTIPLEcast,unnamedcast18883USEDMULTIPLEcast,unnamedcast18881USEDMULTIPLEcast,unnamedcast18879USEDMULTIPLEcast,unnamedcast18877USEDMULTIPLEcast,({inp[407:400]}),unnamedcast18873USEDMULTIPLEcast,unnamedcast18871USEDMULTIPLEcast,unnamedcast18869USEDMULTIPLEcast,unnamedcast18867USEDMULTIPLEcast,unnamedcast18865USEDMULTIPLEcast,unnamedcast18863USEDMULTIPLEcast,unnamedcast18861USEDMULTIPLEcast,unnamedcast18859USEDMULTIPLEcast,unnamedcast18857USEDMULTIPLEcast,unnamedcast18855USEDMULTIPLEcast,unnamedcast18853USEDMULTIPLEcast,unnamedcast18851USEDMULTIPLEcast,unnamedcast18849USEDMULTIPLEcast,unnamedcast18847USEDMULTIPLEcast,unnamedcast18845USEDMULTIPLEcast,({inp[271:264]}),unnamedcast18841USEDMULTIPLEcast,unnamedcast18839USEDMULTIPLEcast,unnamedcast18837USEDMULTIPLEcast,unnamedcast18835USEDMULTIPLEcast,unnamedcast18833USEDMULTIPLEcast,unnamedcast18831USEDMULTIPLEcast,unnamedcast18829USEDMULTIPLEcast,unnamedcast18827USEDMULTIPLEcast,unnamedcast18825USEDMULTIPLEcast,unnamedcast18823USEDMULTIPLEcast,unnamedcast18821USEDMULTIPLEcast,unnamedcast18819USEDMULTIPLEcast,unnamedcast18817USEDMULTIPLEcast,unnamedcast18815USEDMULTIPLEcast,unnamedcast18813USEDMULTIPLEcast,({inp[135:128]}),unnamedcast18809USEDMULTIPLEcast,unnamedcast18807USEDMULTIPLEcast,unnamedcast18805USEDMULTIPLEcast,unnamedcast18803USEDMULTIPLEcast,unnamedcast18801USEDMULTIPLEcast,unnamedcast18799USEDMULTIPLEcast,unnamedcast18797USEDMULTIPLEcast,unnamedcast18795USEDMULTIPLEcast,unnamedcast18793USEDMULTIPLEcast,unnamedcast18791USEDMULTIPLEcast,unnamedcast18789USEDMULTIPLEcast,unnamedcast18787USEDMULTIPLEcast,unnamedcast18785USEDMULTIPLEcast,unnamedcast18783USEDMULTIPLEcast,unnamedcast18781USEDMULTIPLEcast},{unnamedcast19289USEDMULTIPLEcast,unnamedcast19287USEDMULTIPLEcast,unnamedcast19285USEDMULTIPLEcast,unnamedcast19283USEDMULTIPLEcast,unnamedcast19281USEDMULTIPLEcast,unnamedcast19279USEDMULTIPLEcast,unnamedcast19277USEDMULTIPLEcast,unnamedcast19275USEDMULTIPLEcast,unnamedcast19273USEDMULTIPLEcast,unnamedcast19271USEDMULTIPLEcast,unnamedcast19269USEDMULTIPLEcast,unnamedcast19267USEDMULTIPLEcast,unnamedcast19265USEDMULTIPLEcast,unnamedcast19263USEDMULTIPLEcast,unnamedcast19261USEDMULTIPLEcast,({inp[2047:2040]}),unnamedcast19257USEDMULTIPLEcast,unnamedcast19255USEDMULTIPLEcast,unnamedcast19253USEDMULTIPLEcast,unnamedcast19251USEDMULTIPLEcast,unnamedcast19249USEDMULTIPLEcast,unnamedcast19247USEDMULTIPLEcast,unnamedcast19245USEDMULTIPLEcast,unnamedcast19243USEDMULTIPLEcast,unnamedcast19241USEDMULTIPLEcast,unnamedcast19239USEDMULTIPLEcast,unnamedcast19237USEDMULTIPLEcast,unnamedcast19235USEDMULTIPLEcast,unnamedcast19233USEDMULTIPLEcast,unnamedcast19231USEDMULTIPLEcast,unnamedcast19229USEDMULTIPLEcast,({inp[1911:1904]}),unnamedcast19225USEDMULTIPLEcast,unnamedcast19223USEDMULTIPLEcast,unnamedcast19221USEDMULTIPLEcast,unnamedcast19219USEDMULTIPLEcast,unnamedcast19217USEDMULTIPLEcast,unnamedcast19215USEDMULTIPLEcast,unnamedcast19213USEDMULTIPLEcast,unnamedcast19211USEDMULTIPLEcast,unnamedcast19209USEDMULTIPLEcast,unnamedcast19207USEDMULTIPLEcast,unnamedcast19205USEDMULTIPLEcast,unnamedcast19203USEDMULTIPLEcast,unnamedcast19201USEDMULTIPLEcast,unnamedcast19199USEDMULTIPLEcast,unnamedcast19197USEDMULTIPLEcast,({inp[1775:1768]}),unnamedcast19193USEDMULTIPLEcast,unnamedcast19191USEDMULTIPLEcast,unnamedcast19189USEDMULTIPLEcast,unnamedcast19187USEDMULTIPLEcast,unnamedcast19185USEDMULTIPLEcast,unnamedcast19183USEDMULTIPLEcast,unnamedcast19181USEDMULTIPLEcast,unnamedcast19179USEDMULTIPLEcast,unnamedcast19177USEDMULTIPLEcast,unnamedcast19175USEDMULTIPLEcast,unnamedcast19173USEDMULTIPLEcast,unnamedcast19171USEDMULTIPLEcast,unnamedcast19169USEDMULTIPLEcast,unnamedcast19167USEDMULTIPLEcast,unnamedcast19165USEDMULTIPLEcast,({inp[1639:1632]}),unnamedcast19161USEDMULTIPLEcast,unnamedcast19159USEDMULTIPLEcast,unnamedcast19157USEDMULTIPLEcast,unnamedcast19155USEDMULTIPLEcast,unnamedcast19153USEDMULTIPLEcast,unnamedcast19151USEDMULTIPLEcast,unnamedcast19149USEDMULTIPLEcast,unnamedcast19147USEDMULTIPLEcast,unnamedcast19145USEDMULTIPLEcast,unnamedcast19143USEDMULTIPLEcast,unnamedcast19141USEDMULTIPLEcast,unnamedcast19139USEDMULTIPLEcast,unnamedcast19137USEDMULTIPLEcast,unnamedcast19135USEDMULTIPLEcast,unnamedcast19133USEDMULTIPLEcast,({inp[1503:1496]}),unnamedcast19129USEDMULTIPLEcast,unnamedcast19127USEDMULTIPLEcast,unnamedcast19125USEDMULTIPLEcast,unnamedcast19123USEDMULTIPLEcast,unnamedcast19121USEDMULTIPLEcast,unnamedcast19119USEDMULTIPLEcast,unnamedcast19117USEDMULTIPLEcast,unnamedcast19115USEDMULTIPLEcast,unnamedcast19113USEDMULTIPLEcast,unnamedcast19111USEDMULTIPLEcast,unnamedcast19109USEDMULTIPLEcast,unnamedcast19107USEDMULTIPLEcast,unnamedcast19105USEDMULTIPLEcast,unnamedcast19103USEDMULTIPLEcast,unnamedcast19101USEDMULTIPLEcast,({inp[1367:1360]}),unnamedcast19097USEDMULTIPLEcast,unnamedcast19095USEDMULTIPLEcast,unnamedcast19093USEDMULTIPLEcast,unnamedcast19091USEDMULTIPLEcast,unnamedcast19089USEDMULTIPLEcast,unnamedcast19087USEDMULTIPLEcast,unnamedcast19085USEDMULTIPLEcast,unnamedcast19083USEDMULTIPLEcast,unnamedcast19081USEDMULTIPLEcast,unnamedcast19079USEDMULTIPLEcast,unnamedcast19077USEDMULTIPLEcast,unnamedcast19075USEDMULTIPLEcast,unnamedcast19073USEDMULTIPLEcast,unnamedcast19071USEDMULTIPLEcast,unnamedcast19069USEDMULTIPLEcast,({inp[1231:1224]}),unnamedcast19065USEDMULTIPLEcast,unnamedcast19063USEDMULTIPLEcast,unnamedcast19061USEDMULTIPLEcast,unnamedcast19059USEDMULTIPLEcast,unnamedcast19057USEDMULTIPLEcast,unnamedcast19055USEDMULTIPLEcast,unnamedcast19053USEDMULTIPLEcast,unnamedcast19051USEDMULTIPLEcast,unnamedcast19049USEDMULTIPLEcast,unnamedcast19047USEDMULTIPLEcast,unnamedcast19045USEDMULTIPLEcast,unnamedcast19043USEDMULTIPLEcast,unnamedcast19041USEDMULTIPLEcast,unnamedcast19039USEDMULTIPLEcast,unnamedcast19037USEDMULTIPLEcast,({inp[1095:1088]}),unnamedcast19033USEDMULTIPLEcast,unnamedcast19031USEDMULTIPLEcast,unnamedcast19029USEDMULTIPLEcast,unnamedcast19027USEDMULTIPLEcast,unnamedcast19025USEDMULTIPLEcast,unnamedcast19023USEDMULTIPLEcast,unnamedcast19021USEDMULTIPLEcast,unnamedcast19019USEDMULTIPLEcast,unnamedcast19017USEDMULTIPLEcast,unnamedcast19015USEDMULTIPLEcast,unnamedcast19013USEDMULTIPLEcast,unnamedcast19011USEDMULTIPLEcast,unnamedcast19009USEDMULTIPLEcast,unnamedcast19007USEDMULTIPLEcast,unnamedcast19005USEDMULTIPLEcast,({inp[959:952]}),unnamedcast19001USEDMULTIPLEcast,unnamedcast18999USEDMULTIPLEcast,unnamedcast18997USEDMULTIPLEcast,unnamedcast18995USEDMULTIPLEcast,unnamedcast18993USEDMULTIPLEcast,unnamedcast18991USEDMULTIPLEcast,unnamedcast18989USEDMULTIPLEcast,unnamedcast18987USEDMULTIPLEcast,unnamedcast18985USEDMULTIPLEcast,unnamedcast18983USEDMULTIPLEcast,unnamedcast18981USEDMULTIPLEcast,unnamedcast18979USEDMULTIPLEcast,unnamedcast18977USEDMULTIPLEcast,unnamedcast18975USEDMULTIPLEcast,unnamedcast18973USEDMULTIPLEcast,({inp[823:816]}),unnamedcast18969USEDMULTIPLEcast,unnamedcast18967USEDMULTIPLEcast,unnamedcast18965USEDMULTIPLEcast,unnamedcast18963USEDMULTIPLEcast,unnamedcast18961USEDMULTIPLEcast,unnamedcast18959USEDMULTIPLEcast,unnamedcast18957USEDMULTIPLEcast,unnamedcast18955USEDMULTIPLEcast,unnamedcast18953USEDMULTIPLEcast,unnamedcast18951USEDMULTIPLEcast,unnamedcast18949USEDMULTIPLEcast,unnamedcast18947USEDMULTIPLEcast,unnamedcast18945USEDMULTIPLEcast,unnamedcast18943USEDMULTIPLEcast,unnamedcast18941USEDMULTIPLEcast,({inp[687:680]}),unnamedcast18937USEDMULTIPLEcast,unnamedcast18935USEDMULTIPLEcast,unnamedcast18933USEDMULTIPLEcast,unnamedcast18931USEDMULTIPLEcast,unnamedcast18929USEDMULTIPLEcast,unnamedcast18927USEDMULTIPLEcast,unnamedcast18925USEDMULTIPLEcast,unnamedcast18923USEDMULTIPLEcast,unnamedcast18921USEDMULTIPLEcast,unnamedcast18919USEDMULTIPLEcast,unnamedcast18917USEDMULTIPLEcast,unnamedcast18915USEDMULTIPLEcast,unnamedcast18913USEDMULTIPLEcast,unnamedcast18911USEDMULTIPLEcast,unnamedcast18909USEDMULTIPLEcast,({inp[551:544]}),unnamedcast18905USEDMULTIPLEcast,unnamedcast18903USEDMULTIPLEcast,unnamedcast18901USEDMULTIPLEcast,unnamedcast18899USEDMULTIPLEcast,unnamedcast18897USEDMULTIPLEcast,unnamedcast18895USEDMULTIPLEcast,unnamedcast18893USEDMULTIPLEcast,unnamedcast18891USEDMULTIPLEcast,unnamedcast18889USEDMULTIPLEcast,unnamedcast18887USEDMULTIPLEcast,unnamedcast18885USEDMULTIPLEcast,unnamedcast18883USEDMULTIPLEcast,unnamedcast18881USEDMULTIPLEcast,unnamedcast18879USEDMULTIPLEcast,unnamedcast18877USEDMULTIPLEcast,({inp[415:408]}),unnamedcast18873USEDMULTIPLEcast,unnamedcast18871USEDMULTIPLEcast,unnamedcast18869USEDMULTIPLEcast,unnamedcast18867USEDMULTIPLEcast,unnamedcast18865USEDMULTIPLEcast,unnamedcast18863USEDMULTIPLEcast,unnamedcast18861USEDMULTIPLEcast,unnamedcast18859USEDMULTIPLEcast,unnamedcast18857USEDMULTIPLEcast,unnamedcast18855USEDMULTIPLEcast,unnamedcast18853USEDMULTIPLEcast,unnamedcast18851USEDMULTIPLEcast,unnamedcast18849USEDMULTIPLEcast,unnamedcast18847USEDMULTIPLEcast,unnamedcast18845USEDMULTIPLEcast,({inp[279:272]}),unnamedcast18841USEDMULTIPLEcast,unnamedcast18839USEDMULTIPLEcast,unnamedcast18837USEDMULTIPLEcast,unnamedcast18835USEDMULTIPLEcast,unnamedcast18833USEDMULTIPLEcast,unnamedcast18831USEDMULTIPLEcast,unnamedcast18829USEDMULTIPLEcast,unnamedcast18827USEDMULTIPLEcast,unnamedcast18825USEDMULTIPLEcast,unnamedcast18823USEDMULTIPLEcast,unnamedcast18821USEDMULTIPLEcast,unnamedcast18819USEDMULTIPLEcast,unnamedcast18817USEDMULTIPLEcast,unnamedcast18815USEDMULTIPLEcast,unnamedcast18813USEDMULTIPLEcast,({inp[143:136]}),unnamedcast18809USEDMULTIPLEcast,unnamedcast18807USEDMULTIPLEcast,unnamedcast18805USEDMULTIPLEcast,unnamedcast18803USEDMULTIPLEcast,unnamedcast18801USEDMULTIPLEcast,unnamedcast18799USEDMULTIPLEcast,unnamedcast18797USEDMULTIPLEcast,unnamedcast18795USEDMULTIPLEcast,unnamedcast18793USEDMULTIPLEcast,unnamedcast18791USEDMULTIPLEcast,unnamedcast18789USEDMULTIPLEcast,unnamedcast18787USEDMULTIPLEcast,unnamedcast18785USEDMULTIPLEcast,unnamedcast18783USEDMULTIPLEcast,unnamedcast18781USEDMULTIPLEcast,({inp[7:0]})}};
  // function: process pure=true delay=0
endmodule

module MakeHandshake_unpackStencil_uint8_W16_H16_T2(input CLK, input ready_downstream, output ready, input reset, input [2176:0] process_input, output [4096:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  assign ready = ready_downstream;
  wire unnamedbinop21358USEDMULTIPLEbinop;assign unnamedbinop21358USEDMULTIPLEbinop = {(ready_downstream||reset)}; 
  wire unnamedcast21366USEDMULTIPLEcast;assign unnamedcast21366USEDMULTIPLEcast = (process_input[2176]); 
  wire [4095:0] inner_process_output;
  wire validBitDelay_unpackStencil_uint8_W16_H16_T2_pushPop_out;
  always @(posedge CLK) begin if({(~{(unnamedcast21366USEDMULTIPLEcast===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: MakeHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = {validBitDelay_unpackStencil_uint8_W16_H16_T2_pushPop_out,inner_process_output};
  // function: ready pure=true ONLY WIRE
  // function: reset pure=true ONLY WIRE
  // function: process pure=false ONLY WIRE
  ShiftRegister_0_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_validBitDelay_unpackStencil_uint8_W16_H16_T2"})) validBitDelay_unpackStencil_uint8_W16_H16_T2(.CLK(CLK), .CE(unnamedbinop21358USEDMULTIPLEbinop), .sr_input(unnamedcast21366USEDMULTIPLEcast), .pushPop_out(validBitDelay_unpackStencil_uint8_W16_H16_T2_pushPop_out));
  unpackStencil_uint8_W16_H16_T2 #(.INSTANCE_NAME({INSTANCE_NAME,"_inner"})) inner(.CLK(CLK), .process_CE(unnamedbinop21358USEDMULTIPLEbinop), .inp((process_input[2175:0])), .process_output(inner_process_output));
endmodule

module SSR_W16_H16_T1_Auint8(input CLK, input process_valid, input process_CE, input [127:0] inp, output [2047:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  reg [7:0] SR_x0_y0;
  reg [7:0] SR_x1_y0;
  reg [7:0] SR_x2_y0;
  reg [7:0] SR_x3_y0;
  reg [7:0] SR_x4_y0;
  reg [7:0] SR_x5_y0;
  reg [7:0] SR_x6_y0;
  reg [7:0] SR_x7_y0;
  reg [7:0] SR_x8_y0;
  reg [7:0] SR_x9_y0;
  reg [7:0] SR_x10_y0;
  reg [7:0] SR_x11_y0;
  reg [7:0] SR_x12_y0;
  reg [7:0] SR_x13_y0;
  reg [7:0] SR_x14_y0;
  wire [7:0] unnamedcast21400USEDMULTIPLEcast;assign unnamedcast21400USEDMULTIPLEcast = ({inp[7:0]}); 
  reg [7:0] SR_x0_y1;
  reg [7:0] SR_x1_y1;
  reg [7:0] SR_x2_y1;
  reg [7:0] SR_x3_y1;
  reg [7:0] SR_x4_y1;
  reg [7:0] SR_x5_y1;
  reg [7:0] SR_x6_y1;
  reg [7:0] SR_x7_y1;
  reg [7:0] SR_x8_y1;
  reg [7:0] SR_x9_y1;
  reg [7:0] SR_x10_y1;
  reg [7:0] SR_x11_y1;
  reg [7:0] SR_x12_y1;
  reg [7:0] SR_x13_y1;
  reg [7:0] SR_x14_y1;
  wire [7:0] unnamedcast21448USEDMULTIPLEcast;assign unnamedcast21448USEDMULTIPLEcast = ({inp[15:8]}); 
  reg [7:0] SR_x0_y2;
  reg [7:0] SR_x1_y2;
  reg [7:0] SR_x2_y2;
  reg [7:0] SR_x3_y2;
  reg [7:0] SR_x4_y2;
  reg [7:0] SR_x5_y2;
  reg [7:0] SR_x6_y2;
  reg [7:0] SR_x7_y2;
  reg [7:0] SR_x8_y2;
  reg [7:0] SR_x9_y2;
  reg [7:0] SR_x10_y2;
  reg [7:0] SR_x11_y2;
  reg [7:0] SR_x12_y2;
  reg [7:0] SR_x13_y2;
  reg [7:0] SR_x14_y2;
  wire [7:0] unnamedcast21496USEDMULTIPLEcast;assign unnamedcast21496USEDMULTIPLEcast = ({inp[23:16]}); 
  reg [7:0] SR_x0_y3;
  reg [7:0] SR_x1_y3;
  reg [7:0] SR_x2_y3;
  reg [7:0] SR_x3_y3;
  reg [7:0] SR_x4_y3;
  reg [7:0] SR_x5_y3;
  reg [7:0] SR_x6_y3;
  reg [7:0] SR_x7_y3;
  reg [7:0] SR_x8_y3;
  reg [7:0] SR_x9_y3;
  reg [7:0] SR_x10_y3;
  reg [7:0] SR_x11_y3;
  reg [7:0] SR_x12_y3;
  reg [7:0] SR_x13_y3;
  reg [7:0] SR_x14_y3;
  wire [7:0] unnamedcast21544USEDMULTIPLEcast;assign unnamedcast21544USEDMULTIPLEcast = ({inp[31:24]}); 
  reg [7:0] SR_x0_y4;
  reg [7:0] SR_x1_y4;
  reg [7:0] SR_x2_y4;
  reg [7:0] SR_x3_y4;
  reg [7:0] SR_x4_y4;
  reg [7:0] SR_x5_y4;
  reg [7:0] SR_x6_y4;
  reg [7:0] SR_x7_y4;
  reg [7:0] SR_x8_y4;
  reg [7:0] SR_x9_y4;
  reg [7:0] SR_x10_y4;
  reg [7:0] SR_x11_y4;
  reg [7:0] SR_x12_y4;
  reg [7:0] SR_x13_y4;
  reg [7:0] SR_x14_y4;
  wire [7:0] unnamedcast21592USEDMULTIPLEcast;assign unnamedcast21592USEDMULTIPLEcast = ({inp[39:32]}); 
  reg [7:0] SR_x0_y5;
  reg [7:0] SR_x1_y5;
  reg [7:0] SR_x2_y5;
  reg [7:0] SR_x3_y5;
  reg [7:0] SR_x4_y5;
  reg [7:0] SR_x5_y5;
  reg [7:0] SR_x6_y5;
  reg [7:0] SR_x7_y5;
  reg [7:0] SR_x8_y5;
  reg [7:0] SR_x9_y5;
  reg [7:0] SR_x10_y5;
  reg [7:0] SR_x11_y5;
  reg [7:0] SR_x12_y5;
  reg [7:0] SR_x13_y5;
  reg [7:0] SR_x14_y5;
  wire [7:0] unnamedcast21640USEDMULTIPLEcast;assign unnamedcast21640USEDMULTIPLEcast = ({inp[47:40]}); 
  reg [7:0] SR_x0_y6;
  reg [7:0] SR_x1_y6;
  reg [7:0] SR_x2_y6;
  reg [7:0] SR_x3_y6;
  reg [7:0] SR_x4_y6;
  reg [7:0] SR_x5_y6;
  reg [7:0] SR_x6_y6;
  reg [7:0] SR_x7_y6;
  reg [7:0] SR_x8_y6;
  reg [7:0] SR_x9_y6;
  reg [7:0] SR_x10_y6;
  reg [7:0] SR_x11_y6;
  reg [7:0] SR_x12_y6;
  reg [7:0] SR_x13_y6;
  reg [7:0] SR_x14_y6;
  wire [7:0] unnamedcast21688USEDMULTIPLEcast;assign unnamedcast21688USEDMULTIPLEcast = ({inp[55:48]}); 
  reg [7:0] SR_x0_y7;
  reg [7:0] SR_x1_y7;
  reg [7:0] SR_x2_y7;
  reg [7:0] SR_x3_y7;
  reg [7:0] SR_x4_y7;
  reg [7:0] SR_x5_y7;
  reg [7:0] SR_x6_y7;
  reg [7:0] SR_x7_y7;
  reg [7:0] SR_x8_y7;
  reg [7:0] SR_x9_y7;
  reg [7:0] SR_x10_y7;
  reg [7:0] SR_x11_y7;
  reg [7:0] SR_x12_y7;
  reg [7:0] SR_x13_y7;
  reg [7:0] SR_x14_y7;
  wire [7:0] unnamedcast21736USEDMULTIPLEcast;assign unnamedcast21736USEDMULTIPLEcast = ({inp[63:56]}); 
  reg [7:0] SR_x0_y8;
  reg [7:0] SR_x1_y8;
  reg [7:0] SR_x2_y8;
  reg [7:0] SR_x3_y8;
  reg [7:0] SR_x4_y8;
  reg [7:0] SR_x5_y8;
  reg [7:0] SR_x6_y8;
  reg [7:0] SR_x7_y8;
  reg [7:0] SR_x8_y8;
  reg [7:0] SR_x9_y8;
  reg [7:0] SR_x10_y8;
  reg [7:0] SR_x11_y8;
  reg [7:0] SR_x12_y8;
  reg [7:0] SR_x13_y8;
  reg [7:0] SR_x14_y8;
  wire [7:0] unnamedcast21784USEDMULTIPLEcast;assign unnamedcast21784USEDMULTIPLEcast = ({inp[71:64]}); 
  reg [7:0] SR_x0_y9;
  reg [7:0] SR_x1_y9;
  reg [7:0] SR_x2_y9;
  reg [7:0] SR_x3_y9;
  reg [7:0] SR_x4_y9;
  reg [7:0] SR_x5_y9;
  reg [7:0] SR_x6_y9;
  reg [7:0] SR_x7_y9;
  reg [7:0] SR_x8_y9;
  reg [7:0] SR_x9_y9;
  reg [7:0] SR_x10_y9;
  reg [7:0] SR_x11_y9;
  reg [7:0] SR_x12_y9;
  reg [7:0] SR_x13_y9;
  reg [7:0] SR_x14_y9;
  wire [7:0] unnamedcast21832USEDMULTIPLEcast;assign unnamedcast21832USEDMULTIPLEcast = ({inp[79:72]}); 
  reg [7:0] SR_x0_y10;
  reg [7:0] SR_x1_y10;
  reg [7:0] SR_x2_y10;
  reg [7:0] SR_x3_y10;
  reg [7:0] SR_x4_y10;
  reg [7:0] SR_x5_y10;
  reg [7:0] SR_x6_y10;
  reg [7:0] SR_x7_y10;
  reg [7:0] SR_x8_y10;
  reg [7:0] SR_x9_y10;
  reg [7:0] SR_x10_y10;
  reg [7:0] SR_x11_y10;
  reg [7:0] SR_x12_y10;
  reg [7:0] SR_x13_y10;
  reg [7:0] SR_x14_y10;
  wire [7:0] unnamedcast21880USEDMULTIPLEcast;assign unnamedcast21880USEDMULTIPLEcast = ({inp[87:80]}); 
  reg [7:0] SR_x0_y11;
  reg [7:0] SR_x1_y11;
  reg [7:0] SR_x2_y11;
  reg [7:0] SR_x3_y11;
  reg [7:0] SR_x4_y11;
  reg [7:0] SR_x5_y11;
  reg [7:0] SR_x6_y11;
  reg [7:0] SR_x7_y11;
  reg [7:0] SR_x8_y11;
  reg [7:0] SR_x9_y11;
  reg [7:0] SR_x10_y11;
  reg [7:0] SR_x11_y11;
  reg [7:0] SR_x12_y11;
  reg [7:0] SR_x13_y11;
  reg [7:0] SR_x14_y11;
  wire [7:0] unnamedcast21928USEDMULTIPLEcast;assign unnamedcast21928USEDMULTIPLEcast = ({inp[95:88]}); 
  reg [7:0] SR_x0_y12;
  reg [7:0] SR_x1_y12;
  reg [7:0] SR_x2_y12;
  reg [7:0] SR_x3_y12;
  reg [7:0] SR_x4_y12;
  reg [7:0] SR_x5_y12;
  reg [7:0] SR_x6_y12;
  reg [7:0] SR_x7_y12;
  reg [7:0] SR_x8_y12;
  reg [7:0] SR_x9_y12;
  reg [7:0] SR_x10_y12;
  reg [7:0] SR_x11_y12;
  reg [7:0] SR_x12_y12;
  reg [7:0] SR_x13_y12;
  reg [7:0] SR_x14_y12;
  wire [7:0] unnamedcast21976USEDMULTIPLEcast;assign unnamedcast21976USEDMULTIPLEcast = ({inp[103:96]}); 
  reg [7:0] SR_x0_y13;
  reg [7:0] SR_x1_y13;
  reg [7:0] SR_x2_y13;
  reg [7:0] SR_x3_y13;
  reg [7:0] SR_x4_y13;
  reg [7:0] SR_x5_y13;
  reg [7:0] SR_x6_y13;
  reg [7:0] SR_x7_y13;
  reg [7:0] SR_x8_y13;
  reg [7:0] SR_x9_y13;
  reg [7:0] SR_x10_y13;
  reg [7:0] SR_x11_y13;
  reg [7:0] SR_x12_y13;
  reg [7:0] SR_x13_y13;
  reg [7:0] SR_x14_y13;
  wire [7:0] unnamedcast22024USEDMULTIPLEcast;assign unnamedcast22024USEDMULTIPLEcast = ({inp[111:104]}); 
  reg [7:0] SR_x0_y14;
  reg [7:0] SR_x1_y14;
  reg [7:0] SR_x2_y14;
  reg [7:0] SR_x3_y14;
  reg [7:0] SR_x4_y14;
  reg [7:0] SR_x5_y14;
  reg [7:0] SR_x6_y14;
  reg [7:0] SR_x7_y14;
  reg [7:0] SR_x8_y14;
  reg [7:0] SR_x9_y14;
  reg [7:0] SR_x10_y14;
  reg [7:0] SR_x11_y14;
  reg [7:0] SR_x12_y14;
  reg [7:0] SR_x13_y14;
  reg [7:0] SR_x14_y14;
  wire [7:0] unnamedcast22072USEDMULTIPLEcast;assign unnamedcast22072USEDMULTIPLEcast = ({inp[119:112]}); 
  reg [7:0] SR_x0_y15;
  reg [7:0] SR_x1_y15;
  reg [7:0] SR_x2_y15;
  reg [7:0] SR_x3_y15;
  reg [7:0] SR_x4_y15;
  reg [7:0] SR_x5_y15;
  reg [7:0] SR_x6_y15;
  reg [7:0] SR_x7_y15;
  reg [7:0] SR_x8_y15;
  reg [7:0] SR_x9_y15;
  reg [7:0] SR_x10_y15;
  reg [7:0] SR_x11_y15;
  reg [7:0] SR_x12_y15;
  reg [7:0] SR_x13_y15;
  reg [7:0] SR_x14_y15;
  wire [7:0] unnamedcast22120USEDMULTIPLEcast;assign unnamedcast22120USEDMULTIPLEcast = ({inp[127:120]}); 
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x14_y0 <= unnamedcast21400USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x13_y0 <= SR_x14_y0; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x12_y0 <= SR_x13_y0; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x11_y0 <= SR_x12_y0; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x10_y0 <= SR_x11_y0; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x9_y0 <= SR_x10_y0; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x8_y0 <= SR_x9_y0; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x7_y0 <= SR_x8_y0; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x6_y0 <= SR_x7_y0; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x5_y0 <= SR_x6_y0; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x4_y0 <= SR_x5_y0; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x3_y0 <= SR_x4_y0; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x2_y0 <= SR_x3_y0; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x1_y0 <= SR_x2_y0; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x0_y0 <= SR_x1_y0; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x14_y1 <= unnamedcast21448USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x13_y1 <= SR_x14_y1; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x12_y1 <= SR_x13_y1; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x11_y1 <= SR_x12_y1; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x10_y1 <= SR_x11_y1; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x9_y1 <= SR_x10_y1; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x8_y1 <= SR_x9_y1; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x7_y1 <= SR_x8_y1; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x6_y1 <= SR_x7_y1; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x5_y1 <= SR_x6_y1; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x4_y1 <= SR_x5_y1; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x3_y1 <= SR_x4_y1; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x2_y1 <= SR_x3_y1; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x1_y1 <= SR_x2_y1; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x0_y1 <= SR_x1_y1; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x14_y2 <= unnamedcast21496USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x13_y2 <= SR_x14_y2; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x12_y2 <= SR_x13_y2; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x11_y2 <= SR_x12_y2; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x10_y2 <= SR_x11_y2; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x9_y2 <= SR_x10_y2; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x8_y2 <= SR_x9_y2; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x7_y2 <= SR_x8_y2; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x6_y2 <= SR_x7_y2; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x5_y2 <= SR_x6_y2; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x4_y2 <= SR_x5_y2; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x3_y2 <= SR_x4_y2; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x2_y2 <= SR_x3_y2; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x1_y2 <= SR_x2_y2; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x0_y2 <= SR_x1_y2; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x14_y3 <= unnamedcast21544USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x13_y3 <= SR_x14_y3; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x12_y3 <= SR_x13_y3; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x11_y3 <= SR_x12_y3; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x10_y3 <= SR_x11_y3; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x9_y3 <= SR_x10_y3; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x8_y3 <= SR_x9_y3; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x7_y3 <= SR_x8_y3; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x6_y3 <= SR_x7_y3; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x5_y3 <= SR_x6_y3; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x4_y3 <= SR_x5_y3; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x3_y3 <= SR_x4_y3; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x2_y3 <= SR_x3_y3; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x1_y3 <= SR_x2_y3; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x0_y3 <= SR_x1_y3; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x14_y4 <= unnamedcast21592USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x13_y4 <= SR_x14_y4; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x12_y4 <= SR_x13_y4; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x11_y4 <= SR_x12_y4; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x10_y4 <= SR_x11_y4; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x9_y4 <= SR_x10_y4; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x8_y4 <= SR_x9_y4; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x7_y4 <= SR_x8_y4; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x6_y4 <= SR_x7_y4; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x5_y4 <= SR_x6_y4; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x4_y4 <= SR_x5_y4; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x3_y4 <= SR_x4_y4; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x2_y4 <= SR_x3_y4; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x1_y4 <= SR_x2_y4; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x0_y4 <= SR_x1_y4; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x14_y5 <= unnamedcast21640USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x13_y5 <= SR_x14_y5; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x12_y5 <= SR_x13_y5; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x11_y5 <= SR_x12_y5; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x10_y5 <= SR_x11_y5; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x9_y5 <= SR_x10_y5; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x8_y5 <= SR_x9_y5; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x7_y5 <= SR_x8_y5; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x6_y5 <= SR_x7_y5; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x5_y5 <= SR_x6_y5; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x4_y5 <= SR_x5_y5; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x3_y5 <= SR_x4_y5; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x2_y5 <= SR_x3_y5; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x1_y5 <= SR_x2_y5; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x0_y5 <= SR_x1_y5; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x14_y6 <= unnamedcast21688USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x13_y6 <= SR_x14_y6; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x12_y6 <= SR_x13_y6; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x11_y6 <= SR_x12_y6; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x10_y6 <= SR_x11_y6; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x9_y6 <= SR_x10_y6; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x8_y6 <= SR_x9_y6; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x7_y6 <= SR_x8_y6; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x6_y6 <= SR_x7_y6; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x5_y6 <= SR_x6_y6; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x4_y6 <= SR_x5_y6; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x3_y6 <= SR_x4_y6; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x2_y6 <= SR_x3_y6; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x1_y6 <= SR_x2_y6; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x0_y6 <= SR_x1_y6; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x14_y7 <= unnamedcast21736USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x13_y7 <= SR_x14_y7; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x12_y7 <= SR_x13_y7; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x11_y7 <= SR_x12_y7; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x10_y7 <= SR_x11_y7; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x9_y7 <= SR_x10_y7; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x8_y7 <= SR_x9_y7; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x7_y7 <= SR_x8_y7; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x6_y7 <= SR_x7_y7; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x5_y7 <= SR_x6_y7; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x4_y7 <= SR_x5_y7; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x3_y7 <= SR_x4_y7; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x2_y7 <= SR_x3_y7; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x1_y7 <= SR_x2_y7; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x0_y7 <= SR_x1_y7; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x14_y8 <= unnamedcast21784USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x13_y8 <= SR_x14_y8; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x12_y8 <= SR_x13_y8; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x11_y8 <= SR_x12_y8; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x10_y8 <= SR_x11_y8; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x9_y8 <= SR_x10_y8; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x8_y8 <= SR_x9_y8; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x7_y8 <= SR_x8_y8; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x6_y8 <= SR_x7_y8; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x5_y8 <= SR_x6_y8; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x4_y8 <= SR_x5_y8; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x3_y8 <= SR_x4_y8; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x2_y8 <= SR_x3_y8; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x1_y8 <= SR_x2_y8; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x0_y8 <= SR_x1_y8; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x14_y9 <= unnamedcast21832USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x13_y9 <= SR_x14_y9; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x12_y9 <= SR_x13_y9; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x11_y9 <= SR_x12_y9; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x10_y9 <= SR_x11_y9; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x9_y9 <= SR_x10_y9; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x8_y9 <= SR_x9_y9; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x7_y9 <= SR_x8_y9; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x6_y9 <= SR_x7_y9; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x5_y9 <= SR_x6_y9; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x4_y9 <= SR_x5_y9; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x3_y9 <= SR_x4_y9; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x2_y9 <= SR_x3_y9; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x1_y9 <= SR_x2_y9; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x0_y9 <= SR_x1_y9; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x14_y10 <= unnamedcast21880USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x13_y10 <= SR_x14_y10; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x12_y10 <= SR_x13_y10; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x11_y10 <= SR_x12_y10; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x10_y10 <= SR_x11_y10; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x9_y10 <= SR_x10_y10; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x8_y10 <= SR_x9_y10; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x7_y10 <= SR_x8_y10; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x6_y10 <= SR_x7_y10; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x5_y10 <= SR_x6_y10; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x4_y10 <= SR_x5_y10; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x3_y10 <= SR_x4_y10; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x2_y10 <= SR_x3_y10; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x1_y10 <= SR_x2_y10; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x0_y10 <= SR_x1_y10; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x14_y11 <= unnamedcast21928USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x13_y11 <= SR_x14_y11; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x12_y11 <= SR_x13_y11; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x11_y11 <= SR_x12_y11; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x10_y11 <= SR_x11_y11; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x9_y11 <= SR_x10_y11; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x8_y11 <= SR_x9_y11; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x7_y11 <= SR_x8_y11; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x6_y11 <= SR_x7_y11; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x5_y11 <= SR_x6_y11; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x4_y11 <= SR_x5_y11; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x3_y11 <= SR_x4_y11; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x2_y11 <= SR_x3_y11; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x1_y11 <= SR_x2_y11; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x0_y11 <= SR_x1_y11; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x14_y12 <= unnamedcast21976USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x13_y12 <= SR_x14_y12; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x12_y12 <= SR_x13_y12; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x11_y12 <= SR_x12_y12; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x10_y12 <= SR_x11_y12; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x9_y12 <= SR_x10_y12; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x8_y12 <= SR_x9_y12; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x7_y12 <= SR_x8_y12; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x6_y12 <= SR_x7_y12; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x5_y12 <= SR_x6_y12; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x4_y12 <= SR_x5_y12; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x3_y12 <= SR_x4_y12; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x2_y12 <= SR_x3_y12; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x1_y12 <= SR_x2_y12; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x0_y12 <= SR_x1_y12; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x14_y13 <= unnamedcast22024USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x13_y13 <= SR_x14_y13; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x12_y13 <= SR_x13_y13; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x11_y13 <= SR_x12_y13; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x10_y13 <= SR_x11_y13; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x9_y13 <= SR_x10_y13; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x8_y13 <= SR_x9_y13; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x7_y13 <= SR_x8_y13; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x6_y13 <= SR_x7_y13; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x5_y13 <= SR_x6_y13; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x4_y13 <= SR_x5_y13; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x3_y13 <= SR_x4_y13; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x2_y13 <= SR_x3_y13; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x1_y13 <= SR_x2_y13; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x0_y13 <= SR_x1_y13; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x14_y14 <= unnamedcast22072USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x13_y14 <= SR_x14_y14; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x12_y14 <= SR_x13_y14; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x11_y14 <= SR_x12_y14; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x10_y14 <= SR_x11_y14; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x9_y14 <= SR_x10_y14; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x8_y14 <= SR_x9_y14; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x7_y14 <= SR_x8_y14; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x6_y14 <= SR_x7_y14; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x5_y14 <= SR_x6_y14; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x4_y14 <= SR_x5_y14; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x3_y14 <= SR_x4_y14; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x2_y14 <= SR_x3_y14; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x1_y14 <= SR_x2_y14; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x0_y14 <= SR_x1_y14; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x14_y15 <= unnamedcast22120USEDMULTIPLEcast; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x13_y15 <= SR_x14_y15; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x12_y15 <= SR_x13_y15; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x11_y15 <= SR_x12_y15; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x10_y15 <= SR_x11_y15; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x9_y15 <= SR_x10_y15; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x8_y15 <= SR_x9_y15; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x7_y15 <= SR_x8_y15; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x6_y15 <= SR_x7_y15; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x5_y15 <= SR_x6_y15; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x4_y15 <= SR_x5_y15; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x3_y15 <= SR_x4_y15; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x2_y15 <= SR_x3_y15; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x1_y15 <= SR_x2_y15; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_x0_y15 <= SR_x1_y15; end end
  assign process_output = {unnamedcast22120USEDMULTIPLEcast,SR_x14_y15,SR_x13_y15,SR_x12_y15,SR_x11_y15,SR_x10_y15,SR_x9_y15,SR_x8_y15,SR_x7_y15,SR_x6_y15,SR_x5_y15,SR_x4_y15,SR_x3_y15,SR_x2_y15,SR_x1_y15,SR_x0_y15,unnamedcast22072USEDMULTIPLEcast,SR_x14_y14,SR_x13_y14,SR_x12_y14,SR_x11_y14,SR_x10_y14,SR_x9_y14,SR_x8_y14,SR_x7_y14,SR_x6_y14,SR_x5_y14,SR_x4_y14,SR_x3_y14,SR_x2_y14,SR_x1_y14,SR_x0_y14,unnamedcast22024USEDMULTIPLEcast,SR_x14_y13,SR_x13_y13,SR_x12_y13,SR_x11_y13,SR_x10_y13,SR_x9_y13,SR_x8_y13,SR_x7_y13,SR_x6_y13,SR_x5_y13,SR_x4_y13,SR_x3_y13,SR_x2_y13,SR_x1_y13,SR_x0_y13,unnamedcast21976USEDMULTIPLEcast,SR_x14_y12,SR_x13_y12,SR_x12_y12,SR_x11_y12,SR_x10_y12,SR_x9_y12,SR_x8_y12,SR_x7_y12,SR_x6_y12,SR_x5_y12,SR_x4_y12,SR_x3_y12,SR_x2_y12,SR_x1_y12,SR_x0_y12,unnamedcast21928USEDMULTIPLEcast,SR_x14_y11,SR_x13_y11,SR_x12_y11,SR_x11_y11,SR_x10_y11,SR_x9_y11,SR_x8_y11,SR_x7_y11,SR_x6_y11,SR_x5_y11,SR_x4_y11,SR_x3_y11,SR_x2_y11,SR_x1_y11,SR_x0_y11,unnamedcast21880USEDMULTIPLEcast,SR_x14_y10,SR_x13_y10,SR_x12_y10,SR_x11_y10,SR_x10_y10,SR_x9_y10,SR_x8_y10,SR_x7_y10,SR_x6_y10,SR_x5_y10,SR_x4_y10,SR_x3_y10,SR_x2_y10,SR_x1_y10,SR_x0_y10,unnamedcast21832USEDMULTIPLEcast,SR_x14_y9,SR_x13_y9,SR_x12_y9,SR_x11_y9,SR_x10_y9,SR_x9_y9,SR_x8_y9,SR_x7_y9,SR_x6_y9,SR_x5_y9,SR_x4_y9,SR_x3_y9,SR_x2_y9,SR_x1_y9,SR_x0_y9,unnamedcast21784USEDMULTIPLEcast,SR_x14_y8,SR_x13_y8,SR_x12_y8,SR_x11_y8,SR_x10_y8,SR_x9_y8,SR_x8_y8,SR_x7_y8,SR_x6_y8,SR_x5_y8,SR_x4_y8,SR_x3_y8,SR_x2_y8,SR_x1_y8,SR_x0_y8,unnamedcast21736USEDMULTIPLEcast,SR_x14_y7,SR_x13_y7,SR_x12_y7,SR_x11_y7,SR_x10_y7,SR_x9_y7,SR_x8_y7,SR_x7_y7,SR_x6_y7,SR_x5_y7,SR_x4_y7,SR_x3_y7,SR_x2_y7,SR_x1_y7,SR_x0_y7,unnamedcast21688USEDMULTIPLEcast,SR_x14_y6,SR_x13_y6,SR_x12_y6,SR_x11_y6,SR_x10_y6,SR_x9_y6,SR_x8_y6,SR_x7_y6,SR_x6_y6,SR_x5_y6,SR_x4_y6,SR_x3_y6,SR_x2_y6,SR_x1_y6,SR_x0_y6,unnamedcast21640USEDMULTIPLEcast,SR_x14_y5,SR_x13_y5,SR_x12_y5,SR_x11_y5,SR_x10_y5,SR_x9_y5,SR_x8_y5,SR_x7_y5,SR_x6_y5,SR_x5_y5,SR_x4_y5,SR_x3_y5,SR_x2_y5,SR_x1_y5,SR_x0_y5,unnamedcast21592USEDMULTIPLEcast,SR_x14_y4,SR_x13_y4,SR_x12_y4,SR_x11_y4,SR_x10_y4,SR_x9_y4,SR_x8_y4,SR_x7_y4,SR_x6_y4,SR_x5_y4,SR_x4_y4,SR_x3_y4,SR_x2_y4,SR_x1_y4,SR_x0_y4,unnamedcast21544USEDMULTIPLEcast,SR_x14_y3,SR_x13_y3,SR_x12_y3,SR_x11_y3,SR_x10_y3,SR_x9_y3,SR_x8_y3,SR_x7_y3,SR_x6_y3,SR_x5_y3,SR_x4_y3,SR_x3_y3,SR_x2_y3,SR_x1_y3,SR_x0_y3,unnamedcast21496USEDMULTIPLEcast,SR_x14_y2,SR_x13_y2,SR_x12_y2,SR_x11_y2,SR_x10_y2,SR_x9_y2,SR_x8_y2,SR_x7_y2,SR_x6_y2,SR_x5_y2,SR_x4_y2,SR_x3_y2,SR_x2_y2,SR_x1_y2,SR_x0_y2,unnamedcast21448USEDMULTIPLEcast,SR_x14_y1,SR_x13_y1,SR_x12_y1,SR_x11_y1,SR_x10_y1,SR_x9_y1,SR_x8_y1,SR_x7_y1,SR_x6_y1,SR_x5_y1,SR_x4_y1,SR_x3_y1,SR_x2_y1,SR_x1_y1,SR_x0_y1,unnamedcast21400USEDMULTIPLEcast,SR_x14_y0,SR_x13_y0,SR_x12_y0,SR_x11_y0,SR_x10_y0,SR_x9_y0,SR_x8_y0,SR_x7_y0,SR_x6_y0,SR_x5_y0,SR_x4_y0,SR_x3_y0,SR_x2_y0,SR_x1_y0,SR_x0_y0};
  // function: process pure=false delay=0
  // function: reset pure=true delay=0
endmodule

module stencilLinebuffer_Auint8_w831_h495_xmin15_ymin15(input CLK, input process_valid, input CE, input [7:0] process_input, output [2047:0] process_output, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  wire [127:0] stencilLinebuffer_Auint8_w831_h495_xmin15_ymin15_g_process_output;
  reg process_valid_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay1_validunnamednull0_CECE <= process_valid; end end
  reg process_valid_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay2_validunnamednull0_CECE <= process_valid_delay1_validunnamednull0_CECE; end end
  reg process_valid_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay3_validunnamednull0_CECE <= process_valid_delay2_validunnamednull0_CECE; end end
  reg process_valid_delay4_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay4_validunnamednull0_CECE <= process_valid_delay3_validunnamednull0_CECE; end end
  reg process_valid_delay5_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay5_validunnamednull0_CECE <= process_valid_delay4_validunnamednull0_CECE; end end
  reg process_valid_delay6_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay6_validunnamednull0_CECE <= process_valid_delay5_validunnamednull0_CECE; end end
  reg process_valid_delay7_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay7_validunnamednull0_CECE <= process_valid_delay6_validunnamednull0_CECE; end end
  reg process_valid_delay8_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay8_validunnamednull0_CECE <= process_valid_delay7_validunnamednull0_CECE; end end
  reg process_valid_delay9_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay9_validunnamednull0_CECE <= process_valid_delay8_validunnamednull0_CECE; end end
  reg process_valid_delay10_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay10_validunnamednull0_CECE <= process_valid_delay9_validunnamednull0_CECE; end end
  reg process_valid_delay11_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay11_validunnamednull0_CECE <= process_valid_delay10_validunnamednull0_CECE; end end
  reg process_valid_delay12_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay12_validunnamednull0_CECE <= process_valid_delay11_validunnamednull0_CECE; end end
  reg process_valid_delay13_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay13_validunnamednull0_CECE <= process_valid_delay12_validunnamednull0_CECE; end end
  reg process_valid_delay14_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay14_validunnamednull0_CECE <= process_valid_delay13_validunnamednull0_CECE; end end
  reg process_valid_delay15_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay15_validunnamednull0_CECE <= process_valid_delay14_validunnamednull0_CECE; end end
  wire [2047:0] stencilLinebuffer_Auint8_w831_h495_xmin15_ymin15_f_process_output;
  assign process_output = stencilLinebuffer_Auint8_w831_h495_xmin15_ymin15_f_process_output;
  // function: process pure=false delay=15
  // function: reset pure=false delay=0
  linebuffer_w831_h495_T1_ymin_15_Auint8 #(.INSTANCE_NAME({INSTANCE_NAME,"_stencilLinebuffer_Auint8_w831_h495_xmin15_ymin15_g"})) stencilLinebuffer_Auint8_w831_h495_xmin15_ymin15_g(.CLK(CLK), .process_valid(process_valid), .CE(CE), .process_input(process_input), .process_output(stencilLinebuffer_Auint8_w831_h495_xmin15_ymin15_g_process_output), .reset(reset));
  SSR_W16_H16_T1_Auint8 #(.INSTANCE_NAME({INSTANCE_NAME,"_stencilLinebuffer_Auint8_w831_h495_xmin15_ymin15_f"})) stencilLinebuffer_Auint8_w831_h495_xmin15_ymin15_f(.CLK(CLK), .process_valid(process_valid_delay15_validunnamednull0_CECE), .process_CE(CE), .inp(stencilLinebuffer_Auint8_w831_h495_xmin15_ymin15_g_process_output), .process_output(stencilLinebuffer_Auint8_w831_h495_xmin15_ymin15_f_process_output));
endmodule

module MakeHandshake_stencilLinebuffer_Auint8_w831_h495_xmin15_ymin15(input CLK, input ready_downstream, output ready, input reset, input [8:0] process_input, output [2048:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  assign ready = ready_downstream;
  wire unnamedbinop23718USEDMULTIPLEbinop;assign unnamedbinop23718USEDMULTIPLEbinop = {(ready_downstream||reset)}; 
  wire unnamedcast23726USEDMULTIPLEcast;assign unnamedcast23726USEDMULTIPLEcast = (process_input[8]); 
  wire [2047:0] inner_process_output;
  wire validBitDelay_stencilLinebuffer_Auint8_w831_h495_xmin15_ymin15_pushPop_out;
  always @(posedge CLK) begin if({(~{(unnamedcast23726USEDMULTIPLEcast===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: MakeHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = {validBitDelay_stencilLinebuffer_Auint8_w831_h495_xmin15_ymin15_pushPop_out,inner_process_output};
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  ShiftRegister_15_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_validBitDelay_stencilLinebuffer_Auint8_w831_h495_xmin15_ymin15"})) validBitDelay_stencilLinebuffer_Auint8_w831_h495_xmin15_ymin15(.CLK(CLK), .pushPop_valid({(~reset)}), .CE(unnamedbinop23718USEDMULTIPLEbinop), .sr_input(unnamedcast23726USEDMULTIPLEcast), .pushPop_out(validBitDelay_stencilLinebuffer_Auint8_w831_h495_xmin15_ymin15_pushPop_out), .reset(reset));
  stencilLinebuffer_Auint8_w831_h495_xmin15_ymin15 #(.INSTANCE_NAME({INSTANCE_NAME,"_inner"})) inner(.CLK(CLK), .process_valid(unnamedcast23726USEDMULTIPLEcast), .CE(unnamedbinop23718USEDMULTIPLEbinop), .process_input((process_input[7:0])), .process_output(inner_process_output), .reset(reset));
endmodule

module arrayop_uint8_16_16__W1_Hnil(input CLK, input CE, input [2047:0] process_input, output [2047:0] process_output);
parameter INSTANCE_NAME="INST";
  assign process_output = {process_input};
  // function: process pure=true delay=0
  // function: reset pure=true delay=0
endmodule

module MakeHandshake_arrayop_uint8_16_16__W1_Hnil(input CLK, input ready_downstream, output ready, input reset, input [2048:0] process_input, output [2048:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  assign ready = ready_downstream;
  wire unnamedbinop23745USEDMULTIPLEbinop;assign unnamedbinop23745USEDMULTIPLEbinop = {(ready_downstream||reset)}; 
  wire unnamedcast23753USEDMULTIPLEcast;assign unnamedcast23753USEDMULTIPLEcast = (process_input[2048]); 
  wire [2047:0] inner_process_output;
  wire validBitDelay_arrayop_uint8_16_16__W1_Hnil_pushPop_out;
  always @(posedge CLK) begin if({(~{(unnamedcast23753USEDMULTIPLEcast===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: MakeHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = {validBitDelay_arrayop_uint8_16_16__W1_Hnil_pushPop_out,inner_process_output};
  // function: ready pure=true ONLY WIRE
  // function: reset pure=true ONLY WIRE
  // function: process pure=false ONLY WIRE
  ShiftRegister_0_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_validBitDelay_arrayop_uint8_16_16__W1_Hnil"})) validBitDelay_arrayop_uint8_16_16__W1_Hnil(.CLK(CLK), .CE(unnamedbinop23745USEDMULTIPLEbinop), .sr_input(unnamedcast23753USEDMULTIPLEcast), .pushPop_out(validBitDelay_arrayop_uint8_16_16__W1_Hnil_pushPop_out));
  arrayop_uint8_16_16__W1_Hnil #(.INSTANCE_NAME({INSTANCE_NAME,"_inner"})) inner(.CLK(CLK), .CE(unnamedbinop23745USEDMULTIPLEbinop), .process_input((process_input[2047:0])), .process_output(inner_process_output));
endmodule

module sumwrap_uint8_to7(input CLK, input CE, input [15:0] process_input, output [7:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [7:0] unnamedcast23758USEDMULTIPLEcast;assign unnamedcast23758USEDMULTIPLEcast = (process_input[7:0]); 
  assign process_output = (({(unnamedcast23758USEDMULTIPLEcast==(8'd7))})?((8'd0)):({(unnamedcast23758USEDMULTIPLEcast+(process_input[15:8]))}));
  // function: process pure=true delay=0
endmodule

module RegBy_sumwrap_uint8_to7_CEtrue_initnil(input CLK, input set_valid, input CE, input [7:0] set_inp, input setby_valid, input [7:0] setby_inp, output [7:0] SETBY_OUTPUT, output [7:0] GET_OUTPUT);
parameter INSTANCE_NAME="INST";
  reg [7:0] R;
  wire [7:0] regby_inner_process_output;
  always @(posedge CLK) begin if(set_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(setby_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,set_valid})+({4'b0,setby_valid})) > 5'd1) begin $display("error, function 'set' on instance 'R' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [8:0] unnamedcallArbitrate23798USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate23798USEDMULTIPLEcallArbitrate = {(set_valid||setby_valid),((set_valid)?(set_inp):(regby_inner_process_output))}; 
    always @ (posedge CLK) begin if ((unnamedcallArbitrate23798USEDMULTIPLEcallArbitrate[8]) && CE) begin R <= (unnamedcallArbitrate23798USEDMULTIPLEcallArbitrate[7:0]); end end
  assign SETBY_OUTPUT = regby_inner_process_output;
  assign GET_OUTPUT = R;
  // function: set pure=false ONLY WIRE
  // function: setby pure=false ONLY WIRE
  // function: get pure=true ONLY WIRE
  sumwrap_uint8_to7 #(.INSTANCE_NAME({INSTANCE_NAME,"_regby_inner"})) regby_inner(.CLK(CLK), .CE(CE), .process_input({setby_inp,R}), .process_output(regby_inner_process_output));
endmodule

module UpsampleXSeq(input CLK, output ready, input reset, input CE, input process_valid, input [2047:0] inp, output [2048:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  wire [7:0] phase_GET_OUTPUT;
  wire unnamedbinop23807USEDMULTIPLEbinop;assign unnamedbinop23807USEDMULTIPLEbinop = {(phase_GET_OUTPUT==(8'd0))}; 
  assign ready = unnamedbinop23807USEDMULTIPLEbinop;
  reg [2047:0] buffer;
  reg [2047:0] unnamedselect23809_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedselect23809_delay1_validunnamednull0_CECE <= ((unnamedbinop23807USEDMULTIPLEbinop)?(inp):(buffer)); end end
    always @ (posedge CLK) begin if ({(unnamedbinop23807USEDMULTIPLEbinop&&process_valid)} && CE) begin buffer <= inp; end end
  wire [7:0] phase_SETBY_OUTPUT;
  assign process_output = {(1'd1),unnamedselect23809_delay1_validunnamednull0_CECE};
  // function: ready pure=true delay=0
  // function: reset pure=false delay=0
  // function: process pure=false delay=1
  RegBy_sumwrap_uint8_to7_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_phase"})) phase(.CLK(CLK), .set_valid(reset), .CE(CE), .set_inp((8'd0)), .setby_valid(process_valid), .setby_inp((8'd1)), .SETBY_OUTPUT(phase_SETBY_OUTPUT), .GET_OUTPUT(phase_GET_OUTPUT));
endmodule

module WaitOnInput_UpsampleXSeq(input CLK, output ready, input reset, input CE, input process_valid, input [2048:0] process_input, output [2048:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  wire WaitOnInput_inner_ready;
  assign ready = WaitOnInput_inner_ready;
  wire unnamedbinop23875USEDMULTIPLEbinop;assign unnamedbinop23875USEDMULTIPLEbinop = {({({(~WaitOnInput_inner_ready)}||(process_input[2048]))}&&process_valid)}; 
  wire [2048:0] WaitOnInput_inner_process_output;
  reg unnamedbinop23875_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedbinop23875_delay1_validunnamednull0_CECE <= unnamedbinop23875USEDMULTIPLEbinop; end end
  assign process_output = {{((WaitOnInput_inner_process_output[2048])&&unnamedbinop23875_delay1_validunnamednull0_CECE)},(WaitOnInput_inner_process_output[2047:0])};
  // function: ready pure=true delay=0
  // function: reset pure=false delay=0
  // function: process pure=false delay=1
  UpsampleXSeq #(.INSTANCE_NAME({INSTANCE_NAME,"_WaitOnInput_inner"})) WaitOnInput_inner(.CLK(CLK), .ready(WaitOnInput_inner_ready), .reset(reset), .CE(CE), .process_valid(unnamedbinop23875USEDMULTIPLEbinop), .inp((process_input[2047:0])), .process_output(WaitOnInput_inner_process_output));
endmodule

module LiftHandshake_WaitOnInput_UpsampleXSeq(input CLK, input ready_downstream, output ready, input reset, input [2048:0] process_input, output [2048:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire inner_WaitOnInput_UpsampleXSeq_ready;
  assign ready = {(inner_WaitOnInput_UpsampleXSeq_ready&&ready_downstream)};
  wire unnamedbinop23910USEDMULTIPLEbinop;assign unnamedbinop23910USEDMULTIPLEbinop = {(reset||ready_downstream)}; 
  wire unnamedunary23911USEDMULTIPLEunary;assign unnamedunary23911USEDMULTIPLEunary = {(~reset)}; 
  wire [2048:0] inner_WaitOnInput_UpsampleXSeq_process_output;
  wire validBitDelay_WaitOnInput_UpsampleXSeq_pushPop_out;
  wire [2048:0] unnamedtuple23921USEDMULTIPLEtuple;assign unnamedtuple23921USEDMULTIPLEtuple = {{((inner_WaitOnInput_UpsampleXSeq_process_output[2048])&&validBitDelay_WaitOnInput_UpsampleXSeq_pushPop_out)},(inner_WaitOnInput_UpsampleXSeq_process_output[2047:0])}; 
  always @(posedge CLK) begin if({(~{((unnamedtuple23921USEDMULTIPLEtuple[2048])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: output valid bit should not be X!",INSTANCE_NAME); end end
  always @(posedge CLK) begin if({(~{((process_input[2048])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = unnamedtuple23921USEDMULTIPLEtuple;
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  WaitOnInput_UpsampleXSeq #(.INSTANCE_NAME({INSTANCE_NAME,"_inner_WaitOnInput_UpsampleXSeq"})) inner_WaitOnInput_UpsampleXSeq(.CLK(CLK), .ready(inner_WaitOnInput_UpsampleXSeq_ready), .reset(reset), .CE(unnamedbinop23910USEDMULTIPLEbinop), .process_valid(unnamedunary23911USEDMULTIPLEunary), .process_input(process_input), .process_output(inner_WaitOnInput_UpsampleXSeq_process_output));
  ShiftRegister_1_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_validBitDelay_WaitOnInput_UpsampleXSeq"})) validBitDelay_WaitOnInput_UpsampleXSeq(.CLK(CLK), .pushPop_valid(unnamedunary23911USEDMULTIPLEunary), .CE(unnamedbinop23910USEDMULTIPLEbinop), .sr_input((1'd1)), .pushPop_out(validBitDelay_WaitOnInput_UpsampleXSeq_pushPop_out), .reset(reset));
endmodule

module slice_typeuint8_16_16__1_1__xl0_xh0_yl0_yh0(input CLK, input process_CE, input [2047:0] inp, output [2047:0] process_output);
parameter INSTANCE_NAME="INST";
  assign process_output = ({inp[2047:0]});
  // function: process pure=true delay=0
endmodule

module MakeHandshake_slice_typeuint8_16_16__1_1__xl0_xh0_yl0_yh0(input CLK, input ready_downstream, output ready, input reset, input [2048:0] process_input, output [2048:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  assign ready = ready_downstream;
  wire unnamedbinop23955USEDMULTIPLEbinop;assign unnamedbinop23955USEDMULTIPLEbinop = {(ready_downstream||reset)}; 
  wire unnamedcast23963USEDMULTIPLEcast;assign unnamedcast23963USEDMULTIPLEcast = (process_input[2048]); 
  wire [2047:0] inner_process_output;
  wire validBitDelay_slice_typeuint8_16_16__1_1__xl0_xh0_yl0_yh0_pushPop_out;
  always @(posedge CLK) begin if({(~{(unnamedcast23963USEDMULTIPLEcast===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: MakeHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = {validBitDelay_slice_typeuint8_16_16__1_1__xl0_xh0_yl0_yh0_pushPop_out,inner_process_output};
  // function: ready pure=true ONLY WIRE
  // function: reset pure=true ONLY WIRE
  // function: process pure=false ONLY WIRE
  ShiftRegister_0_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_validBitDelay_slice_typeuint8_16_16__1_1__xl0_xh0_yl0_yh0"})) validBitDelay_slice_typeuint8_16_16__1_1__xl0_xh0_yl0_yh0(.CLK(CLK), .CE(unnamedbinop23955USEDMULTIPLEbinop), .sr_input(unnamedcast23963USEDMULTIPLEcast), .pushPop_out(validBitDelay_slice_typeuint8_16_16__1_1__xl0_xh0_yl0_yh0_pushPop_out));
  slice_typeuint8_16_16__1_1__xl0_xh0_yl0_yh0 #(.INSTANCE_NAME({INSTANCE_NAME,"_inner"})) inner(.CLK(CLK), .process_CE(unnamedbinop23955USEDMULTIPLEbinop), .inp((process_input[2047:0])), .process_output(inner_process_output));
endmodule

module Broadcast_2(input CLK, input process_CE, input [2047:0] inp, output [4095:0] process_output);
parameter INSTANCE_NAME="INST";
  assign process_output = {inp,inp};
  // function: process pure=true delay=0
endmodule

module MakeHandshake_Broadcast_2(input CLK, input ready_downstream, output ready, input reset, input [2048:0] process_input, output [4096:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  assign ready = ready_downstream;
  wire unnamedbinop23981USEDMULTIPLEbinop;assign unnamedbinop23981USEDMULTIPLEbinop = {(ready_downstream||reset)}; 
  wire unnamedcast23989USEDMULTIPLEcast;assign unnamedcast23989USEDMULTIPLEcast = (process_input[2048]); 
  wire [4095:0] inner_process_output;
  wire validBitDelay_Broadcast_2_pushPop_out;
  always @(posedge CLK) begin if({(~{(unnamedcast23989USEDMULTIPLEcast===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: MakeHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = {validBitDelay_Broadcast_2_pushPop_out,inner_process_output};
  // function: ready pure=true ONLY WIRE
  // function: reset pure=true ONLY WIRE
  // function: process pure=false ONLY WIRE
  ShiftRegister_0_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_validBitDelay_Broadcast_2"})) validBitDelay_Broadcast_2(.CLK(CLK), .CE(unnamedbinop23981USEDMULTIPLEbinop), .sr_input(unnamedcast23989USEDMULTIPLEcast), .pushPop_out(validBitDelay_Broadcast_2_pushPop_out));
  Broadcast_2 #(.INSTANCE_NAME({INSTANCE_NAME,"_inner"})) inner(.CLK(CLK), .process_CE(unnamedbinop23981USEDMULTIPLEbinop), .inp((process_input[2047:0])), .process_output(inner_process_output));
endmodule

module packTuple_table__0x4782d2f8(input CLK, input ready_downstream, output [1:0] ready, input [8193:0] process_input, output [8192:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [4096:0] unnamedcast24067USEDMULTIPLEcast;assign unnamedcast24067USEDMULTIPLEcast = (process_input[4096:0]); 
  wire unnamedcast24069USEDMULTIPLEcast;assign unnamedcast24069USEDMULTIPLEcast = (unnamedcast24067USEDMULTIPLEcast[4096]); 
  wire [4096:0] unnamedcast24071USEDMULTIPLEcast;assign unnamedcast24071USEDMULTIPLEcast = (process_input[8193:4097]); 
  wire unnamedcast24073USEDMULTIPLEcast;assign unnamedcast24073USEDMULTIPLEcast = (unnamedcast24071USEDMULTIPLEcast[4096]); 
  wire unnamedbinop24082USEDMULTIPLEbinop;assign unnamedbinop24082USEDMULTIPLEbinop = {(unnamedcast24069USEDMULTIPLEcast&&unnamedcast24073USEDMULTIPLEcast)}; 
  wire unnamedbinop24087USEDMULTIPLEbinop;assign unnamedbinop24087USEDMULTIPLEbinop = {(ready_downstream&&unnamedbinop24082USEDMULTIPLEbinop)}; 
  assign ready = {{(unnamedbinop24087USEDMULTIPLEbinop||{(~unnamedcast24073USEDMULTIPLEcast)})},{(unnamedbinop24087USEDMULTIPLEbinop||{(~unnamedcast24069USEDMULTIPLEcast)})}};
  assign process_output = {unnamedbinop24082USEDMULTIPLEbinop,{(unnamedcast24071USEDMULTIPLEcast[4095:0]),(unnamedcast24067USEDMULTIPLEcast[4095:0])}};
  // function: ready pure=true ONLY WIRE
  // function: reset pure=true ONLY WIRE
  // function: process pure=true ONLY WIRE
endmodule

module packTupleArrays_table__0x42b86538(input CLK, input process_CE, input [8191:0] process_input, output [8191:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [4095:0] unnamedcast23994USEDMULTIPLEcast;assign unnamedcast23994USEDMULTIPLEcast = (process_input[4095:0]); 
  wire [4095:0] unnamedcast23998USEDMULTIPLEcast;assign unnamedcast23998USEDMULTIPLEcast = (process_input[8191:4096]); 
  assign process_output = {{({unnamedcast23998USEDMULTIPLEcast[4095:2048]}),({unnamedcast23994USEDMULTIPLEcast[4095:2048]})},{({unnamedcast23998USEDMULTIPLEcast[2047:0]}),({unnamedcast23994USEDMULTIPLEcast[2047:0]})}};
  // function: process pure=true delay=0
endmodule

module MakeHandshake_packTupleArrays_table__0x42b86538(input CLK, input ready_downstream, output ready, input reset, input [8192:0] process_input, output [8192:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  assign ready = ready_downstream;
  wire unnamedbinop24045USEDMULTIPLEbinop;assign unnamedbinop24045USEDMULTIPLEbinop = {(ready_downstream||reset)}; 
  wire unnamedcast24053USEDMULTIPLEcast;assign unnamedcast24053USEDMULTIPLEcast = (process_input[8192]); 
  wire [8191:0] inner_process_output;
  wire validBitDelay_packTupleArrays_table__0x42b86538_pushPop_out;
  always @(posedge CLK) begin if({(~{(unnamedcast24053USEDMULTIPLEcast===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: MakeHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = {validBitDelay_packTupleArrays_table__0x42b86538_pushPop_out,inner_process_output};
  // function: ready pure=true ONLY WIRE
  // function: reset pure=true ONLY WIRE
  // function: process pure=false ONLY WIRE
  ShiftRegister_0_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_validBitDelay_packTupleArrays_table__0x42b86538"})) validBitDelay_packTupleArrays_table__0x42b86538(.CLK(CLK), .CE(unnamedbinop24045USEDMULTIPLEbinop), .sr_input(unnamedcast24053USEDMULTIPLEcast), .pushPop_out(validBitDelay_packTupleArrays_table__0x42b86538_pushPop_out));
  packTupleArrays_table__0x42b86538 #(.INSTANCE_NAME({INSTANCE_NAME,"_inner"})) inner(.CLK(CLK), .process_CE(unnamedbinop24045USEDMULTIPLEbinop), .process_input((process_input[8191:0])), .process_output(inner_process_output));
endmodule

module SoAtoAoSHandshake_W2_H1_table__0x42b86538(input CLK, input ready_downstream, output [1:0] ready, input reset, input [8193:0] process_input, output [8192:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire SoAtoAoSHandshake_W2_H1_table__0x42b86538_f_ready;
  wire [1:0] SoAtoAoSHandshake_W2_H1_table__0x42b86538_g_ready;
  assign ready = SoAtoAoSHandshake_W2_H1_table__0x42b86538_g_ready;
  wire [8192:0] SoAtoAoSHandshake_W2_H1_table__0x42b86538_g_process_output;
  wire [8192:0] SoAtoAoSHandshake_W2_H1_table__0x42b86538_f_process_output;
  assign process_output = SoAtoAoSHandshake_W2_H1_table__0x42b86538_f_process_output;
  // function: ready pure=true ONLY WIRE
  // function: reset pure=true ONLY WIRE
  // function: process pure=false ONLY WIRE
  packTuple_table__0x4782d2f8 #(.INSTANCE_NAME({INSTANCE_NAME,"_SoAtoAoSHandshake_W2_H1_table__0x42b86538_g"})) SoAtoAoSHandshake_W2_H1_table__0x42b86538_g(.CLK(CLK), .ready_downstream(SoAtoAoSHandshake_W2_H1_table__0x42b86538_f_ready), .ready(SoAtoAoSHandshake_W2_H1_table__0x42b86538_g_ready), .process_input(process_input), .process_output(SoAtoAoSHandshake_W2_H1_table__0x42b86538_g_process_output));
  MakeHandshake_packTupleArrays_table__0x42b86538 #(.INSTANCE_NAME({INSTANCE_NAME,"_SoAtoAoSHandshake_W2_H1_table__0x42b86538_f"})) SoAtoAoSHandshake_W2_H1_table__0x42b86538_f(.CLK(CLK), .ready_downstream(ready_downstream), .ready(SoAtoAoSHandshake_W2_H1_table__0x42b86538_f_ready), .reset(reset), .process_input(SoAtoAoSHandshake_W2_H1_table__0x42b86538_g_process_output), .process_output(SoAtoAoSHandshake_W2_H1_table__0x42b86538_f_process_output));
endmodule

module packTupleArrays_table__0x4293c570(input CLK, input process_CE, input [4095:0] process_input, output [4095:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [2047:0] unnamedcast24118USEDMULTIPLEcast;assign unnamedcast24118USEDMULTIPLEcast = (process_input[2047:0]); 
  wire [2047:0] unnamedcast24122USEDMULTIPLEcast;assign unnamedcast24122USEDMULTIPLEcast = (process_input[4095:2048]); 
  assign process_output = {{({unnamedcast24122USEDMULTIPLEcast[2047:2040]}),({unnamedcast24118USEDMULTIPLEcast[2047:2040]})},{({unnamedcast24122USEDMULTIPLEcast[2039:2032]}),({unnamedcast24118USEDMULTIPLEcast[2039:2032]})},{({unnamedcast24122USEDMULTIPLEcast[2031:2024]}),({unnamedcast24118USEDMULTIPLEcast[2031:2024]})},{({unnamedcast24122USEDMULTIPLEcast[2023:2016]}),({unnamedcast24118USEDMULTIPLEcast[2023:2016]})},{({unnamedcast24122USEDMULTIPLEcast[2015:2008]}),({unnamedcast24118USEDMULTIPLEcast[2015:2008]})},{({unnamedcast24122USEDMULTIPLEcast[2007:2000]}),({unnamedcast24118USEDMULTIPLEcast[2007:2000]})},{({unnamedcast24122USEDMULTIPLEcast[1999:1992]}),({unnamedcast24118USEDMULTIPLEcast[1999:1992]})},{({unnamedcast24122USEDMULTIPLEcast[1991:1984]}),({unnamedcast24118USEDMULTIPLEcast[1991:1984]})},{({unnamedcast24122USEDMULTIPLEcast[1983:1976]}),({unnamedcast24118USEDMULTIPLEcast[1983:1976]})},{({unnamedcast24122USEDMULTIPLEcast[1975:1968]}),({unnamedcast24118USEDMULTIPLEcast[1975:1968]})},{({unnamedcast24122USEDMULTIPLEcast[1967:1960]}),({unnamedcast24118USEDMULTIPLEcast[1967:1960]})},{({unnamedcast24122USEDMULTIPLEcast[1959:1952]}),({unnamedcast24118USEDMULTIPLEcast[1959:1952]})},{({unnamedcast24122USEDMULTIPLEcast[1951:1944]}),({unnamedcast24118USEDMULTIPLEcast[1951:1944]})},{({unnamedcast24122USEDMULTIPLEcast[1943:1936]}),({unnamedcast24118USEDMULTIPLEcast[1943:1936]})},{({unnamedcast24122USEDMULTIPLEcast[1935:1928]}),({unnamedcast24118USEDMULTIPLEcast[1935:1928]})},{({unnamedcast24122USEDMULTIPLEcast[1927:1920]}),({unnamedcast24118USEDMULTIPLEcast[1927:1920]})},{({unnamedcast24122USEDMULTIPLEcast[1919:1912]}),({unnamedcast24118USEDMULTIPLEcast[1919:1912]})},{({unnamedcast24122USEDMULTIPLEcast[1911:1904]}),({unnamedcast24118USEDMULTIPLEcast[1911:1904]})},{({unnamedcast24122USEDMULTIPLEcast[1903:1896]}),({unnamedcast24118USEDMULTIPLEcast[1903:1896]})},{({unnamedcast24122USEDMULTIPLEcast[1895:1888]}),({unnamedcast24118USEDMULTIPLEcast[1895:1888]})},{({unnamedcast24122USEDMULTIPLEcast[1887:1880]}),({unnamedcast24118USEDMULTIPLEcast[1887:1880]})},{({unnamedcast24122USEDMULTIPLEcast[1879:1872]}),({unnamedcast24118USEDMULTIPLEcast[1879:1872]})},{({unnamedcast24122USEDMULTIPLEcast[1871:1864]}),({unnamedcast24118USEDMULTIPLEcast[1871:1864]})},{({unnamedcast24122USEDMULTIPLEcast[1863:1856]}),({unnamedcast24118USEDMULTIPLEcast[1863:1856]})},{({unnamedcast24122USEDMULTIPLEcast[1855:1848]}),({unnamedcast24118USEDMULTIPLEcast[1855:1848]})},{({unnamedcast24122USEDMULTIPLEcast[1847:1840]}),({unnamedcast24118USEDMULTIPLEcast[1847:1840]})},{({unnamedcast24122USEDMULTIPLEcast[1839:1832]}),({unnamedcast24118USEDMULTIPLEcast[1839:1832]})},{({unnamedcast24122USEDMULTIPLEcast[1831:1824]}),({unnamedcast24118USEDMULTIPLEcast[1831:1824]})},{({unnamedcast24122USEDMULTIPLEcast[1823:1816]}),({unnamedcast24118USEDMULTIPLEcast[1823:1816]})},{({unnamedcast24122USEDMULTIPLEcast[1815:1808]}),({unnamedcast24118USEDMULTIPLEcast[1815:1808]})},{({unnamedcast24122USEDMULTIPLEcast[1807:1800]}),({unnamedcast24118USEDMULTIPLEcast[1807:1800]})},{({unnamedcast24122USEDMULTIPLEcast[1799:1792]}),({unnamedcast24118USEDMULTIPLEcast[1799:1792]})},{({unnamedcast24122USEDMULTIPLEcast[1791:1784]}),({unnamedcast24118USEDMULTIPLEcast[1791:1784]})},{({unnamedcast24122USEDMULTIPLEcast[1783:1776]}),({unnamedcast24118USEDMULTIPLEcast[1783:1776]})},{({unnamedcast24122USEDMULTIPLEcast[1775:1768]}),({unnamedcast24118USEDMULTIPLEcast[1775:1768]})},{({unnamedcast24122USEDMULTIPLEcast[1767:1760]}),({unnamedcast24118USEDMULTIPLEcast[1767:1760]})},{({unnamedcast24122USEDMULTIPLEcast[1759:1752]}),({unnamedcast24118USEDMULTIPLEcast[1759:1752]})},{({unnamedcast24122USEDMULTIPLEcast[1751:1744]}),({unnamedcast24118USEDMULTIPLEcast[1751:1744]})},{({unnamedcast24122USEDMULTIPLEcast[1743:1736]}),({unnamedcast24118USEDMULTIPLEcast[1743:1736]})},{({unnamedcast24122USEDMULTIPLEcast[1735:1728]}),({unnamedcast24118USEDMULTIPLEcast[1735:1728]})},{({unnamedcast24122USEDMULTIPLEcast[1727:1720]}),({unnamedcast24118USEDMULTIPLEcast[1727:1720]})},{({unnamedcast24122USEDMULTIPLEcast[1719:1712]}),({unnamedcast24118USEDMULTIPLEcast[1719:1712]})},{({unnamedcast24122USEDMULTIPLEcast[1711:1704]}),({unnamedcast24118USEDMULTIPLEcast[1711:1704]})},{({unnamedcast24122USEDMULTIPLEcast[1703:1696]}),({unnamedcast24118USEDMULTIPLEcast[1703:1696]})},{({unnamedcast24122USEDMULTIPLEcast[1695:1688]}),({unnamedcast24118USEDMULTIPLEcast[1695:1688]})},{({unnamedcast24122USEDMULTIPLEcast[1687:1680]}),({unnamedcast24118USEDMULTIPLEcast[1687:1680]})},{({unnamedcast24122USEDMULTIPLEcast[1679:1672]}),({unnamedcast24118USEDMULTIPLEcast[1679:1672]})},{({unnamedcast24122USEDMULTIPLEcast[1671:1664]}),({unnamedcast24118USEDMULTIPLEcast[1671:1664]})},{({unnamedcast24122USEDMULTIPLEcast[1663:1656]}),({unnamedcast24118USEDMULTIPLEcast[1663:1656]})},{({unnamedcast24122USEDMULTIPLEcast[1655:1648]}),({unnamedcast24118USEDMULTIPLEcast[1655:1648]})},{({unnamedcast24122USEDMULTIPLEcast[1647:1640]}),({unnamedcast24118USEDMULTIPLEcast[1647:1640]})},{({unnamedcast24122USEDMULTIPLEcast[1639:1632]}),({unnamedcast24118USEDMULTIPLEcast[1639:1632]})},{({unnamedcast24122USEDMULTIPLEcast[1631:1624]}),({unnamedcast24118USEDMULTIPLEcast[1631:1624]})},{({unnamedcast24122USEDMULTIPLEcast[1623:1616]}),({unnamedcast24118USEDMULTIPLEcast[1623:1616]})},{({unnamedcast24122USEDMULTIPLEcast[1615:1608]}),({unnamedcast24118USEDMULTIPLEcast[1615:1608]})},{({unnamedcast24122USEDMULTIPLEcast[1607:1600]}),({unnamedcast24118USEDMULTIPLEcast[1607:1600]})},{({unnamedcast24122USEDMULTIPLEcast[1599:1592]}),({unnamedcast24118USEDMULTIPLEcast[1599:1592]})},{({unnamedcast24122USEDMULTIPLEcast[1591:1584]}),({unnamedcast24118USEDMULTIPLEcast[1591:1584]})},{({unnamedcast24122USEDMULTIPLEcast[1583:1576]}),({unnamedcast24118USEDMULTIPLEcast[1583:1576]})},{({unnamedcast24122USEDMULTIPLEcast[1575:1568]}),({unnamedcast24118USEDMULTIPLEcast[1575:1568]})},{({unnamedcast24122USEDMULTIPLEcast[1567:1560]}),({unnamedcast24118USEDMULTIPLEcast[1567:1560]})},{({unnamedcast24122USEDMULTIPLEcast[1559:1552]}),({unnamedcast24118USEDMULTIPLEcast[1559:1552]})},{({unnamedcast24122USEDMULTIPLEcast[1551:1544]}),({unnamedcast24118USEDMULTIPLEcast[1551:1544]})},{({unnamedcast24122USEDMULTIPLEcast[1543:1536]}),({unnamedcast24118USEDMULTIPLEcast[1543:1536]})},{({unnamedcast24122USEDMULTIPLEcast[1535:1528]}),({unnamedcast24118USEDMULTIPLEcast[1535:1528]})},{({unnamedcast24122USEDMULTIPLEcast[1527:1520]}),({unnamedcast24118USEDMULTIPLEcast[1527:1520]})},{({unnamedcast24122USEDMULTIPLEcast[1519:1512]}),({unnamedcast24118USEDMULTIPLEcast[1519:1512]})},{({unnamedcast24122USEDMULTIPLEcast[1511:1504]}),({unnamedcast24118USEDMULTIPLEcast[1511:1504]})},{({unnamedcast24122USEDMULTIPLEcast[1503:1496]}),({unnamedcast24118USEDMULTIPLEcast[1503:1496]})},{({unnamedcast24122USEDMULTIPLEcast[1495:1488]}),({unnamedcast24118USEDMULTIPLEcast[1495:1488]})},{({unnamedcast24122USEDMULTIPLEcast[1487:1480]}),({unnamedcast24118USEDMULTIPLEcast[1487:1480]})},{({unnamedcast24122USEDMULTIPLEcast[1479:1472]}),({unnamedcast24118USEDMULTIPLEcast[1479:1472]})},{({unnamedcast24122USEDMULTIPLEcast[1471:1464]}),({unnamedcast24118USEDMULTIPLEcast[1471:1464]})},{({unnamedcast24122USEDMULTIPLEcast[1463:1456]}),({unnamedcast24118USEDMULTIPLEcast[1463:1456]})},{({unnamedcast24122USEDMULTIPLEcast[1455:1448]}),({unnamedcast24118USEDMULTIPLEcast[1455:1448]})},{({unnamedcast24122USEDMULTIPLEcast[1447:1440]}),({unnamedcast24118USEDMULTIPLEcast[1447:1440]})},{({unnamedcast24122USEDMULTIPLEcast[1439:1432]}),({unnamedcast24118USEDMULTIPLEcast[1439:1432]})},{({unnamedcast24122USEDMULTIPLEcast[1431:1424]}),({unnamedcast24118USEDMULTIPLEcast[1431:1424]})},{({unnamedcast24122USEDMULTIPLEcast[1423:1416]}),({unnamedcast24118USEDMULTIPLEcast[1423:1416]})},{({unnamedcast24122USEDMULTIPLEcast[1415:1408]}),({unnamedcast24118USEDMULTIPLEcast[1415:1408]})},{({unnamedcast24122USEDMULTIPLEcast[1407:1400]}),({unnamedcast24118USEDMULTIPLEcast[1407:1400]})},{({unnamedcast24122USEDMULTIPLEcast[1399:1392]}),({unnamedcast24118USEDMULTIPLEcast[1399:1392]})},{({unnamedcast24122USEDMULTIPLEcast[1391:1384]}),({unnamedcast24118USEDMULTIPLEcast[1391:1384]})},{({unnamedcast24122USEDMULTIPLEcast[1383:1376]}),({unnamedcast24118USEDMULTIPLEcast[1383:1376]})},{({unnamedcast24122USEDMULTIPLEcast[1375:1368]}),({unnamedcast24118USEDMULTIPLEcast[1375:1368]})},{({unnamedcast24122USEDMULTIPLEcast[1367:1360]}),({unnamedcast24118USEDMULTIPLEcast[1367:1360]})},{({unnamedcast24122USEDMULTIPLEcast[1359:1352]}),({unnamedcast24118USEDMULTIPLEcast[1359:1352]})},{({unnamedcast24122USEDMULTIPLEcast[1351:1344]}),({unnamedcast24118USEDMULTIPLEcast[1351:1344]})},{({unnamedcast24122USEDMULTIPLEcast[1343:1336]}),({unnamedcast24118USEDMULTIPLEcast[1343:1336]})},{({unnamedcast24122USEDMULTIPLEcast[1335:1328]}),({unnamedcast24118USEDMULTIPLEcast[1335:1328]})},{({unnamedcast24122USEDMULTIPLEcast[1327:1320]}),({unnamedcast24118USEDMULTIPLEcast[1327:1320]})},{({unnamedcast24122USEDMULTIPLEcast[1319:1312]}),({unnamedcast24118USEDMULTIPLEcast[1319:1312]})},{({unnamedcast24122USEDMULTIPLEcast[1311:1304]}),({unnamedcast24118USEDMULTIPLEcast[1311:1304]})},{({unnamedcast24122USEDMULTIPLEcast[1303:1296]}),({unnamedcast24118USEDMULTIPLEcast[1303:1296]})},{({unnamedcast24122USEDMULTIPLEcast[1295:1288]}),({unnamedcast24118USEDMULTIPLEcast[1295:1288]})},{({unnamedcast24122USEDMULTIPLEcast[1287:1280]}),({unnamedcast24118USEDMULTIPLEcast[1287:1280]})},{({unnamedcast24122USEDMULTIPLEcast[1279:1272]}),({unnamedcast24118USEDMULTIPLEcast[1279:1272]})},{({unnamedcast24122USEDMULTIPLEcast[1271:1264]}),({unnamedcast24118USEDMULTIPLEcast[1271:1264]})},{({unnamedcast24122USEDMULTIPLEcast[1263:1256]}),({unnamedcast24118USEDMULTIPLEcast[1263:1256]})},{({unnamedcast24122USEDMULTIPLEcast[1255:1248]}),({unnamedcast24118USEDMULTIPLEcast[1255:1248]})},{({unnamedcast24122USEDMULTIPLEcast[1247:1240]}),({unnamedcast24118USEDMULTIPLEcast[1247:1240]})},{({unnamedcast24122USEDMULTIPLEcast[1239:1232]}),({unnamedcast24118USEDMULTIPLEcast[1239:1232]})},{({unnamedcast24122USEDMULTIPLEcast[1231:1224]}),({unnamedcast24118USEDMULTIPLEcast[1231:1224]})},{({unnamedcast24122USEDMULTIPLEcast[1223:1216]}),({unnamedcast24118USEDMULTIPLEcast[1223:1216]})},{({unnamedcast24122USEDMULTIPLEcast[1215:1208]}),({unnamedcast24118USEDMULTIPLEcast[1215:1208]})},{({unnamedcast24122USEDMULTIPLEcast[1207:1200]}),({unnamedcast24118USEDMULTIPLEcast[1207:1200]})},{({unnamedcast24122USEDMULTIPLEcast[1199:1192]}),({unnamedcast24118USEDMULTIPLEcast[1199:1192]})},{({unnamedcast24122USEDMULTIPLEcast[1191:1184]}),({unnamedcast24118USEDMULTIPLEcast[1191:1184]})},{({unnamedcast24122USEDMULTIPLEcast[1183:1176]}),({unnamedcast24118USEDMULTIPLEcast[1183:1176]})},{({unnamedcast24122USEDMULTIPLEcast[1175:1168]}),({unnamedcast24118USEDMULTIPLEcast[1175:1168]})},{({unnamedcast24122USEDMULTIPLEcast[1167:1160]}),({unnamedcast24118USEDMULTIPLEcast[1167:1160]})},{({unnamedcast24122USEDMULTIPLEcast[1159:1152]}),({unnamedcast24118USEDMULTIPLEcast[1159:1152]})},{({unnamedcast24122USEDMULTIPLEcast[1151:1144]}),({unnamedcast24118USEDMULTIPLEcast[1151:1144]})},{({unnamedcast24122USEDMULTIPLEcast[1143:1136]}),({unnamedcast24118USEDMULTIPLEcast[1143:1136]})},{({unnamedcast24122USEDMULTIPLEcast[1135:1128]}),({unnamedcast24118USEDMULTIPLEcast[1135:1128]})},{({unnamedcast24122USEDMULTIPLEcast[1127:1120]}),({unnamedcast24118USEDMULTIPLEcast[1127:1120]})},{({unnamedcast24122USEDMULTIPLEcast[1119:1112]}),({unnamedcast24118USEDMULTIPLEcast[1119:1112]})},{({unnamedcast24122USEDMULTIPLEcast[1111:1104]}),({unnamedcast24118USEDMULTIPLEcast[1111:1104]})},{({unnamedcast24122USEDMULTIPLEcast[1103:1096]}),({unnamedcast24118USEDMULTIPLEcast[1103:1096]})},{({unnamedcast24122USEDMULTIPLEcast[1095:1088]}),({unnamedcast24118USEDMULTIPLEcast[1095:1088]})},{({unnamedcast24122USEDMULTIPLEcast[1087:1080]}),({unnamedcast24118USEDMULTIPLEcast[1087:1080]})},{({unnamedcast24122USEDMULTIPLEcast[1079:1072]}),({unnamedcast24118USEDMULTIPLEcast[1079:1072]})},{({unnamedcast24122USEDMULTIPLEcast[1071:1064]}),({unnamedcast24118USEDMULTIPLEcast[1071:1064]})},{({unnamedcast24122USEDMULTIPLEcast[1063:1056]}),({unnamedcast24118USEDMULTIPLEcast[1063:1056]})},{({unnamedcast24122USEDMULTIPLEcast[1055:1048]}),({unnamedcast24118USEDMULTIPLEcast[1055:1048]})},{({unnamedcast24122USEDMULTIPLEcast[1047:1040]}),({unnamedcast24118USEDMULTIPLEcast[1047:1040]})},{({unnamedcast24122USEDMULTIPLEcast[1039:1032]}),({unnamedcast24118USEDMULTIPLEcast[1039:1032]})},{({unnamedcast24122USEDMULTIPLEcast[1031:1024]}),({unnamedcast24118USEDMULTIPLEcast[1031:1024]})},{({unnamedcast24122USEDMULTIPLEcast[1023:1016]}),({unnamedcast24118USEDMULTIPLEcast[1023:1016]})},{({unnamedcast24122USEDMULTIPLEcast[1015:1008]}),({unnamedcast24118USEDMULTIPLEcast[1015:1008]})},{({unnamedcast24122USEDMULTIPLEcast[1007:1000]}),({unnamedcast24118USEDMULTIPLEcast[1007:1000]})},{({unnamedcast24122USEDMULTIPLEcast[999:992]}),({unnamedcast24118USEDMULTIPLEcast[999:992]})},{({unnamedcast24122USEDMULTIPLEcast[991:984]}),({unnamedcast24118USEDMULTIPLEcast[991:984]})},{({unnamedcast24122USEDMULTIPLEcast[983:976]}),({unnamedcast24118USEDMULTIPLEcast[983:976]})},{({unnamedcast24122USEDMULTIPLEcast[975:968]}),({unnamedcast24118USEDMULTIPLEcast[975:968]})},{({unnamedcast24122USEDMULTIPLEcast[967:960]}),({unnamedcast24118USEDMULTIPLEcast[967:960]})},{({unnamedcast24122USEDMULTIPLEcast[959:952]}),({unnamedcast24118USEDMULTIPLEcast[959:952]})},{({unnamedcast24122USEDMULTIPLEcast[951:944]}),({unnamedcast24118USEDMULTIPLEcast[951:944]})},{({unnamedcast24122USEDMULTIPLEcast[943:936]}),({unnamedcast24118USEDMULTIPLEcast[943:936]})},{({unnamedcast24122USEDMULTIPLEcast[935:928]}),({unnamedcast24118USEDMULTIPLEcast[935:928]})},{({unnamedcast24122USEDMULTIPLEcast[927:920]}),({unnamedcast24118USEDMULTIPLEcast[927:920]})},{({unnamedcast24122USEDMULTIPLEcast[919:912]}),({unnamedcast24118USEDMULTIPLEcast[919:912]})},{({unnamedcast24122USEDMULTIPLEcast[911:904]}),({unnamedcast24118USEDMULTIPLEcast[911:904]})},{({unnamedcast24122USEDMULTIPLEcast[903:896]}),({unnamedcast24118USEDMULTIPLEcast[903:896]})},{({unnamedcast24122USEDMULTIPLEcast[895:888]}),({unnamedcast24118USEDMULTIPLEcast[895:888]})},{({unnamedcast24122USEDMULTIPLEcast[887:880]}),({unnamedcast24118USEDMULTIPLEcast[887:880]})},{({unnamedcast24122USEDMULTIPLEcast[879:872]}),({unnamedcast24118USEDMULTIPLEcast[879:872]})},{({unnamedcast24122USEDMULTIPLEcast[871:864]}),({unnamedcast24118USEDMULTIPLEcast[871:864]})},{({unnamedcast24122USEDMULTIPLEcast[863:856]}),({unnamedcast24118USEDMULTIPLEcast[863:856]})},{({unnamedcast24122USEDMULTIPLEcast[855:848]}),({unnamedcast24118USEDMULTIPLEcast[855:848]})},{({unnamedcast24122USEDMULTIPLEcast[847:840]}),({unnamedcast24118USEDMULTIPLEcast[847:840]})},{({unnamedcast24122USEDMULTIPLEcast[839:832]}),({unnamedcast24118USEDMULTIPLEcast[839:832]})},{({unnamedcast24122USEDMULTIPLEcast[831:824]}),({unnamedcast24118USEDMULTIPLEcast[831:824]})},{({unnamedcast24122USEDMULTIPLEcast[823:816]}),({unnamedcast24118USEDMULTIPLEcast[823:816]})},{({unnamedcast24122USEDMULTIPLEcast[815:808]}),({unnamedcast24118USEDMULTIPLEcast[815:808]})},{({unnamedcast24122USEDMULTIPLEcast[807:800]}),({unnamedcast24118USEDMULTIPLEcast[807:800]})},{({unnamedcast24122USEDMULTIPLEcast[799:792]}),({unnamedcast24118USEDMULTIPLEcast[799:792]})},{({unnamedcast24122USEDMULTIPLEcast[791:784]}),({unnamedcast24118USEDMULTIPLEcast[791:784]})},{({unnamedcast24122USEDMULTIPLEcast[783:776]}),({unnamedcast24118USEDMULTIPLEcast[783:776]})},{({unnamedcast24122USEDMULTIPLEcast[775:768]}),({unnamedcast24118USEDMULTIPLEcast[775:768]})},{({unnamedcast24122USEDMULTIPLEcast[767:760]}),({unnamedcast24118USEDMULTIPLEcast[767:760]})},{({unnamedcast24122USEDMULTIPLEcast[759:752]}),({unnamedcast24118USEDMULTIPLEcast[759:752]})},{({unnamedcast24122USEDMULTIPLEcast[751:744]}),({unnamedcast24118USEDMULTIPLEcast[751:744]})},{({unnamedcast24122USEDMULTIPLEcast[743:736]}),({unnamedcast24118USEDMULTIPLEcast[743:736]})},{({unnamedcast24122USEDMULTIPLEcast[735:728]}),({unnamedcast24118USEDMULTIPLEcast[735:728]})},{({unnamedcast24122USEDMULTIPLEcast[727:720]}),({unnamedcast24118USEDMULTIPLEcast[727:720]})},{({unnamedcast24122USEDMULTIPLEcast[719:712]}),({unnamedcast24118USEDMULTIPLEcast[719:712]})},{({unnamedcast24122USEDMULTIPLEcast[711:704]}),({unnamedcast24118USEDMULTIPLEcast[711:704]})},{({unnamedcast24122USEDMULTIPLEcast[703:696]}),({unnamedcast24118USEDMULTIPLEcast[703:696]})},{({unnamedcast24122USEDMULTIPLEcast[695:688]}),({unnamedcast24118USEDMULTIPLEcast[695:688]})},{({unnamedcast24122USEDMULTIPLEcast[687:680]}),({unnamedcast24118USEDMULTIPLEcast[687:680]})},{({unnamedcast24122USEDMULTIPLEcast[679:672]}),({unnamedcast24118USEDMULTIPLEcast[679:672]})},{({unnamedcast24122USEDMULTIPLEcast[671:664]}),({unnamedcast24118USEDMULTIPLEcast[671:664]})},{({unnamedcast24122USEDMULTIPLEcast[663:656]}),({unnamedcast24118USEDMULTIPLEcast[663:656]})},{({unnamedcast24122USEDMULTIPLEcast[655:648]}),({unnamedcast24118USEDMULTIPLEcast[655:648]})},{({unnamedcast24122USEDMULTIPLEcast[647:640]}),({unnamedcast24118USEDMULTIPLEcast[647:640]})},{({unnamedcast24122USEDMULTIPLEcast[639:632]}),({unnamedcast24118USEDMULTIPLEcast[639:632]})},{({unnamedcast24122USEDMULTIPLEcast[631:624]}),({unnamedcast24118USEDMULTIPLEcast[631:624]})},{({unnamedcast24122USEDMULTIPLEcast[623:616]}),({unnamedcast24118USEDMULTIPLEcast[623:616]})},{({unnamedcast24122USEDMULTIPLEcast[615:608]}),({unnamedcast24118USEDMULTIPLEcast[615:608]})},{({unnamedcast24122USEDMULTIPLEcast[607:600]}),({unnamedcast24118USEDMULTIPLEcast[607:600]})},{({unnamedcast24122USEDMULTIPLEcast[599:592]}),({unnamedcast24118USEDMULTIPLEcast[599:592]})},{({unnamedcast24122USEDMULTIPLEcast[591:584]}),({unnamedcast24118USEDMULTIPLEcast[591:584]})},{({unnamedcast24122USEDMULTIPLEcast[583:576]}),({unnamedcast24118USEDMULTIPLEcast[583:576]})},{({unnamedcast24122USEDMULTIPLEcast[575:568]}),({unnamedcast24118USEDMULTIPLEcast[575:568]})},{({unnamedcast24122USEDMULTIPLEcast[567:560]}),({unnamedcast24118USEDMULTIPLEcast[567:560]})},{({unnamedcast24122USEDMULTIPLEcast[559:552]}),({unnamedcast24118USEDMULTIPLEcast[559:552]})},{({unnamedcast24122USEDMULTIPLEcast[551:544]}),({unnamedcast24118USEDMULTIPLEcast[551:544]})},{({unnamedcast24122USEDMULTIPLEcast[543:536]}),({unnamedcast24118USEDMULTIPLEcast[543:536]})},{({unnamedcast24122USEDMULTIPLEcast[535:528]}),({unnamedcast24118USEDMULTIPLEcast[535:528]})},{({unnamedcast24122USEDMULTIPLEcast[527:520]}),({unnamedcast24118USEDMULTIPLEcast[527:520]})},{({unnamedcast24122USEDMULTIPLEcast[519:512]}),({unnamedcast24118USEDMULTIPLEcast[519:512]})},{({unnamedcast24122USEDMULTIPLEcast[511:504]}),({unnamedcast24118USEDMULTIPLEcast[511:504]})},{({unnamedcast24122USEDMULTIPLEcast[503:496]}),({unnamedcast24118USEDMULTIPLEcast[503:496]})},{({unnamedcast24122USEDMULTIPLEcast[495:488]}),({unnamedcast24118USEDMULTIPLEcast[495:488]})},{({unnamedcast24122USEDMULTIPLEcast[487:480]}),({unnamedcast24118USEDMULTIPLEcast[487:480]})},{({unnamedcast24122USEDMULTIPLEcast[479:472]}),({unnamedcast24118USEDMULTIPLEcast[479:472]})},{({unnamedcast24122USEDMULTIPLEcast[471:464]}),({unnamedcast24118USEDMULTIPLEcast[471:464]})},{({unnamedcast24122USEDMULTIPLEcast[463:456]}),({unnamedcast24118USEDMULTIPLEcast[463:456]})},{({unnamedcast24122USEDMULTIPLEcast[455:448]}),({unnamedcast24118USEDMULTIPLEcast[455:448]})},{({unnamedcast24122USEDMULTIPLEcast[447:440]}),({unnamedcast24118USEDMULTIPLEcast[447:440]})},{({unnamedcast24122USEDMULTIPLEcast[439:432]}),({unnamedcast24118USEDMULTIPLEcast[439:432]})},{({unnamedcast24122USEDMULTIPLEcast[431:424]}),({unnamedcast24118USEDMULTIPLEcast[431:424]})},{({unnamedcast24122USEDMULTIPLEcast[423:416]}),({unnamedcast24118USEDMULTIPLEcast[423:416]})},{({unnamedcast24122USEDMULTIPLEcast[415:408]}),({unnamedcast24118USEDMULTIPLEcast[415:408]})},{({unnamedcast24122USEDMULTIPLEcast[407:400]}),({unnamedcast24118USEDMULTIPLEcast[407:400]})},{({unnamedcast24122USEDMULTIPLEcast[399:392]}),({unnamedcast24118USEDMULTIPLEcast[399:392]})},{({unnamedcast24122USEDMULTIPLEcast[391:384]}),({unnamedcast24118USEDMULTIPLEcast[391:384]})},{({unnamedcast24122USEDMULTIPLEcast[383:376]}),({unnamedcast24118USEDMULTIPLEcast[383:376]})},{({unnamedcast24122USEDMULTIPLEcast[375:368]}),({unnamedcast24118USEDMULTIPLEcast[375:368]})},{({unnamedcast24122USEDMULTIPLEcast[367:360]}),({unnamedcast24118USEDMULTIPLEcast[367:360]})},{({unnamedcast24122USEDMULTIPLEcast[359:352]}),({unnamedcast24118USEDMULTIPLEcast[359:352]})},{({unnamedcast24122USEDMULTIPLEcast[351:344]}),({unnamedcast24118USEDMULTIPLEcast[351:344]})},{({unnamedcast24122USEDMULTIPLEcast[343:336]}),({unnamedcast24118USEDMULTIPLEcast[343:336]})},{({unnamedcast24122USEDMULTIPLEcast[335:328]}),({unnamedcast24118USEDMULTIPLEcast[335:328]})},{({unnamedcast24122USEDMULTIPLEcast[327:320]}),({unnamedcast24118USEDMULTIPLEcast[327:320]})},{({unnamedcast24122USEDMULTIPLEcast[319:312]}),({unnamedcast24118USEDMULTIPLEcast[319:312]})},{({unnamedcast24122USEDMULTIPLEcast[311:304]}),({unnamedcast24118USEDMULTIPLEcast[311:304]})},{({unnamedcast24122USEDMULTIPLEcast[303:296]}),({unnamedcast24118USEDMULTIPLEcast[303:296]})},{({unnamedcast24122USEDMULTIPLEcast[295:288]}),({unnamedcast24118USEDMULTIPLEcast[295:288]})},{({unnamedcast24122USEDMULTIPLEcast[287:280]}),({unnamedcast24118USEDMULTIPLEcast[287:280]})},{({unnamedcast24122USEDMULTIPLEcast[279:272]}),({unnamedcast24118USEDMULTIPLEcast[279:272]})},{({unnamedcast24122USEDMULTIPLEcast[271:264]}),({unnamedcast24118USEDMULTIPLEcast[271:264]})},{({unnamedcast24122USEDMULTIPLEcast[263:256]}),({unnamedcast24118USEDMULTIPLEcast[263:256]})},{({unnamedcast24122USEDMULTIPLEcast[255:248]}),({unnamedcast24118USEDMULTIPLEcast[255:248]})},{({unnamedcast24122USEDMULTIPLEcast[247:240]}),({unnamedcast24118USEDMULTIPLEcast[247:240]})},{({unnamedcast24122USEDMULTIPLEcast[239:232]}),({unnamedcast24118USEDMULTIPLEcast[239:232]})},{({unnamedcast24122USEDMULTIPLEcast[231:224]}),({unnamedcast24118USEDMULTIPLEcast[231:224]})},{({unnamedcast24122USEDMULTIPLEcast[223:216]}),({unnamedcast24118USEDMULTIPLEcast[223:216]})},{({unnamedcast24122USEDMULTIPLEcast[215:208]}),({unnamedcast24118USEDMULTIPLEcast[215:208]})},{({unnamedcast24122USEDMULTIPLEcast[207:200]}),({unnamedcast24118USEDMULTIPLEcast[207:200]})},{({unnamedcast24122USEDMULTIPLEcast[199:192]}),({unnamedcast24118USEDMULTIPLEcast[199:192]})},{({unnamedcast24122USEDMULTIPLEcast[191:184]}),({unnamedcast24118USEDMULTIPLEcast[191:184]})},{({unnamedcast24122USEDMULTIPLEcast[183:176]}),({unnamedcast24118USEDMULTIPLEcast[183:176]})},{({unnamedcast24122USEDMULTIPLEcast[175:168]}),({unnamedcast24118USEDMULTIPLEcast[175:168]})},{({unnamedcast24122USEDMULTIPLEcast[167:160]}),({unnamedcast24118USEDMULTIPLEcast[167:160]})},{({unnamedcast24122USEDMULTIPLEcast[159:152]}),({unnamedcast24118USEDMULTIPLEcast[159:152]})},{({unnamedcast24122USEDMULTIPLEcast[151:144]}),({unnamedcast24118USEDMULTIPLEcast[151:144]})},{({unnamedcast24122USEDMULTIPLEcast[143:136]}),({unnamedcast24118USEDMULTIPLEcast[143:136]})},{({unnamedcast24122USEDMULTIPLEcast[135:128]}),({unnamedcast24118USEDMULTIPLEcast[135:128]})},{({unnamedcast24122USEDMULTIPLEcast[127:120]}),({unnamedcast24118USEDMULTIPLEcast[127:120]})},{({unnamedcast24122USEDMULTIPLEcast[119:112]}),({unnamedcast24118USEDMULTIPLEcast[119:112]})},{({unnamedcast24122USEDMULTIPLEcast[111:104]}),({unnamedcast24118USEDMULTIPLEcast[111:104]})},{({unnamedcast24122USEDMULTIPLEcast[103:96]}),({unnamedcast24118USEDMULTIPLEcast[103:96]})},{({unnamedcast24122USEDMULTIPLEcast[95:88]}),({unnamedcast24118USEDMULTIPLEcast[95:88]})},{({unnamedcast24122USEDMULTIPLEcast[87:80]}),({unnamedcast24118USEDMULTIPLEcast[87:80]})},{({unnamedcast24122USEDMULTIPLEcast[79:72]}),({unnamedcast24118USEDMULTIPLEcast[79:72]})},{({unnamedcast24122USEDMULTIPLEcast[71:64]}),({unnamedcast24118USEDMULTIPLEcast[71:64]})},{({unnamedcast24122USEDMULTIPLEcast[63:56]}),({unnamedcast24118USEDMULTIPLEcast[63:56]})},{({unnamedcast24122USEDMULTIPLEcast[55:48]}),({unnamedcast24118USEDMULTIPLEcast[55:48]})},{({unnamedcast24122USEDMULTIPLEcast[47:40]}),({unnamedcast24118USEDMULTIPLEcast[47:40]})},{({unnamedcast24122USEDMULTIPLEcast[39:32]}),({unnamedcast24118USEDMULTIPLEcast[39:32]})},{({unnamedcast24122USEDMULTIPLEcast[31:24]}),({unnamedcast24118USEDMULTIPLEcast[31:24]})},{({unnamedcast24122USEDMULTIPLEcast[23:16]}),({unnamedcast24118USEDMULTIPLEcast[23:16]})},{({unnamedcast24122USEDMULTIPLEcast[15:8]}),({unnamedcast24118USEDMULTIPLEcast[15:8]})},{({unnamedcast24122USEDMULTIPLEcast[7:0]}),({unnamedcast24118USEDMULTIPLEcast[7:0]})}};
  // function: process pure=true delay=0
endmodule

module map_packTupleArrays_table__0x4293c570_W2_H1(input CLK, input process_CE, input [8191:0] process_input, output [8191:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [4095:0] inner0_0_process_output;
  wire [4095:0] inner1_0_process_output;
  assign process_output = {inner1_0_process_output,inner0_0_process_output};
  // function: process pure=true delay=0
  packTupleArrays_table__0x4293c570 #(.INSTANCE_NAME({INSTANCE_NAME,"_inner0_0"})) inner0_0(.CLK(CLK), .process_CE(process_CE), .process_input(({process_input[4095:0]})), .process_output(inner0_0_process_output));
  packTupleArrays_table__0x4293c570 #(.INSTANCE_NAME({INSTANCE_NAME,"_inner1_0"})) inner1_0(.CLK(CLK), .process_CE(process_CE), .process_input(({process_input[8191:4096]})), .process_output(inner1_0_process_output));
endmodule

module MakeHandshake_map_packTupleArrays_table__0x4293c570_W2_H1(input CLK, input ready_downstream, output ready, input reset, input [8192:0] process_input, output [8192:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  assign ready = ready_downstream;
  wire unnamedbinop29273USEDMULTIPLEbinop;assign unnamedbinop29273USEDMULTIPLEbinop = {(ready_downstream||reset)}; 
  wire unnamedcast29281USEDMULTIPLEcast;assign unnamedcast29281USEDMULTIPLEcast = (process_input[8192]); 
  wire [8191:0] inner_process_output;
  wire validBitDelay_map_packTupleArrays_table__0x4293c570_W2_H1_pushPop_out;
  always @(posedge CLK) begin if({(~{(unnamedcast29281USEDMULTIPLEcast===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: MakeHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = {validBitDelay_map_packTupleArrays_table__0x4293c570_W2_H1_pushPop_out,inner_process_output};
  // function: ready pure=true ONLY WIRE
  // function: reset pure=true ONLY WIRE
  // function: process pure=false ONLY WIRE
  ShiftRegister_0_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_validBitDelay_map_packTupleArrays_table__0x4293c570_W2_H1"})) validBitDelay_map_packTupleArrays_table__0x4293c570_W2_H1(.CLK(CLK), .CE(unnamedbinop29273USEDMULTIPLEbinop), .sr_input(unnamedcast29281USEDMULTIPLEcast), .pushPop_out(validBitDelay_map_packTupleArrays_table__0x4293c570_W2_H1_pushPop_out));
  map_packTupleArrays_table__0x4293c570_W2_H1 #(.INSTANCE_NAME({INSTANCE_NAME,"_inner"})) inner(.CLK(CLK), .process_CE(unnamedbinop29273USEDMULTIPLEbinop), .process_input((process_input[8191:0])), .process_output(inner_process_output));
endmodule

module constSeq_table__0x44c9de70_T8(input CLK, input process_valid, input process_CE, output [15:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  reg [15:0] SR_1 = {8'd190,8'd191};
  reg [15:0] SR_2 = {8'd188,8'd189};
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_1 <= SR_2; end end
  reg [15:0] SR_3 = {8'd186,8'd187};
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_2 <= SR_3; end end
  reg [15:0] SR_4 = {8'd184,8'd185};
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_3 <= SR_4; end end
  reg [15:0] SR_5 = {8'd182,8'd183};
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_4 <= SR_5; end end
  reg [15:0] SR_6 = {8'd180,8'd181};
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_5 <= SR_6; end end
  reg [15:0] SR_7 = {8'd178,8'd179};
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_6 <= SR_7; end end
  reg [15:0] SR_8 = {8'd176,8'd177};
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_7 <= SR_8; end end
    always @ (posedge CLK) begin if (process_valid && process_CE) begin SR_8 <= SR_1; end end
  assign process_output = SR_1;
  // function: process pure=false delay=0
  // function: reset pure=true delay=0
endmodule

module absoluteDiff(input CLK, input process_CE, input [15:0] abs_inp, output [15:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [8:0] unnamedcast29319;assign unnamedcast29319 = {1'b0,({abs_inp[7:0]})};  // wire for int size extend (cast)
  wire [8:0] unnamedcast29322;assign unnamedcast29322 = {1'b0,({abs_inp[15:8]})};  // wire for int size extend (cast)
  wire [9:0] unnamedcast29323;assign unnamedcast29323 = { {1{unnamedcast29319[8]}},unnamedcast29319[8:0]}; // wire for $signed
  wire [9:0] unnamedcast29324;assign unnamedcast29324 = { {1{unnamedcast29322[8]}},unnamedcast29322[8:0]}; // wire for $signed
  reg [9:0] unnamedbinop29325_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop29325_delay1_validunnamednull0_CEprocess_CE <= {($signed(unnamedcast29323)-$signed(unnamedcast29324))}; end end
  reg [9:0] unnamedunary29326_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedunary29326_delay1_validunnamednull0_CEprocess_CE <= {((unnamedbinop29325_delay1_validunnamednull0_CEprocess_CE[9])?(-unnamedbinop29325_delay1_validunnamednull0_CEprocess_CE):(unnamedbinop29325_delay1_validunnamednull0_CEprocess_CE))}; end end
  reg [15:0] unnamedcast29330_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast29330_delay1_validunnamednull0_CEprocess_CE <= (16'd0); end end
  reg [15:0] unnamedcast29330_delay2_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast29330_delay2_validunnamednull0_CEprocess_CE <= unnamedcast29330_delay1_validunnamednull0_CEprocess_CE; end end
  reg [15:0] unnamedbinop29331_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop29331_delay1_validunnamednull0_CEprocess_CE <= {({6'b0,unnamedunary29326_delay1_validunnamednull0_CEprocess_CE}<<<unnamedcast29330_delay2_validunnamednull0_CEprocess_CE)}; end end
  assign process_output = {unnamedbinop29331_delay1_validunnamednull0_CEprocess_CE};
  // function: process pure=true delay=3
endmodule

module map_absoluteDiff_W16_H16(input CLK, input process_CE, input [4095:0] process_input, output [4095:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] inner0_0_process_output;
  wire [15:0] inner1_0_process_output;
  wire [15:0] inner2_0_process_output;
  wire [15:0] inner3_0_process_output;
  wire [15:0] inner4_0_process_output;
  wire [15:0] inner5_0_process_output;
  wire [15:0] inner6_0_process_output;
  wire [15:0] inner7_0_process_output;
  wire [15:0] inner8_0_process_output;
  wire [15:0] inner9_0_process_output;
  wire [15:0] inner10_0_process_output;
  wire [15:0] inner11_0_process_output;
  wire [15:0] inner12_0_process_output;
  wire [15:0] inner13_0_process_output;
  wire [15:0] inner14_0_process_output;
  wire [15:0] inner15_0_process_output;
  wire [15:0] inner0_1_process_output;
  wire [15:0] inner1_1_process_output;
  wire [15:0] inner2_1_process_output;
  wire [15:0] inner3_1_process_output;
  wire [15:0] inner4_1_process_output;
  wire [15:0] inner5_1_process_output;
  wire [15:0] inner6_1_process_output;
  wire [15:0] inner7_1_process_output;
  wire [15:0] inner8_1_process_output;
  wire [15:0] inner9_1_process_output;
  wire [15:0] inner10_1_process_output;
  wire [15:0] inner11_1_process_output;
  wire [15:0] inner12_1_process_output;
  wire [15:0] inner13_1_process_output;
  wire [15:0] inner14_1_process_output;
  wire [15:0] inner15_1_process_output;
  wire [15:0] inner0_2_process_output;
  wire [15:0] inner1_2_process_output;
  wire [15:0] inner2_2_process_output;
  wire [15:0] inner3_2_process_output;
  wire [15:0] inner4_2_process_output;
  wire [15:0] inner5_2_process_output;
  wire [15:0] inner6_2_process_output;
  wire [15:0] inner7_2_process_output;
  wire [15:0] inner8_2_process_output;
  wire [15:0] inner9_2_process_output;
  wire [15:0] inner10_2_process_output;
  wire [15:0] inner11_2_process_output;
  wire [15:0] inner12_2_process_output;
  wire [15:0] inner13_2_process_output;
  wire [15:0] inner14_2_process_output;
  wire [15:0] inner15_2_process_output;
  wire [15:0] inner0_3_process_output;
  wire [15:0] inner1_3_process_output;
  wire [15:0] inner2_3_process_output;
  wire [15:0] inner3_3_process_output;
  wire [15:0] inner4_3_process_output;
  wire [15:0] inner5_3_process_output;
  wire [15:0] inner6_3_process_output;
  wire [15:0] inner7_3_process_output;
  wire [15:0] inner8_3_process_output;
  wire [15:0] inner9_3_process_output;
  wire [15:0] inner10_3_process_output;
  wire [15:0] inner11_3_process_output;
  wire [15:0] inner12_3_process_output;
  wire [15:0] inner13_3_process_output;
  wire [15:0] inner14_3_process_output;
  wire [15:0] inner15_3_process_output;
  wire [15:0] inner0_4_process_output;
  wire [15:0] inner1_4_process_output;
  wire [15:0] inner2_4_process_output;
  wire [15:0] inner3_4_process_output;
  wire [15:0] inner4_4_process_output;
  wire [15:0] inner5_4_process_output;
  wire [15:0] inner6_4_process_output;
  wire [15:0] inner7_4_process_output;
  wire [15:0] inner8_4_process_output;
  wire [15:0] inner9_4_process_output;
  wire [15:0] inner10_4_process_output;
  wire [15:0] inner11_4_process_output;
  wire [15:0] inner12_4_process_output;
  wire [15:0] inner13_4_process_output;
  wire [15:0] inner14_4_process_output;
  wire [15:0] inner15_4_process_output;
  wire [15:0] inner0_5_process_output;
  wire [15:0] inner1_5_process_output;
  wire [15:0] inner2_5_process_output;
  wire [15:0] inner3_5_process_output;
  wire [15:0] inner4_5_process_output;
  wire [15:0] inner5_5_process_output;
  wire [15:0] inner6_5_process_output;
  wire [15:0] inner7_5_process_output;
  wire [15:0] inner8_5_process_output;
  wire [15:0] inner9_5_process_output;
  wire [15:0] inner10_5_process_output;
  wire [15:0] inner11_5_process_output;
  wire [15:0] inner12_5_process_output;
  wire [15:0] inner13_5_process_output;
  wire [15:0] inner14_5_process_output;
  wire [15:0] inner15_5_process_output;
  wire [15:0] inner0_6_process_output;
  wire [15:0] inner1_6_process_output;
  wire [15:0] inner2_6_process_output;
  wire [15:0] inner3_6_process_output;
  wire [15:0] inner4_6_process_output;
  wire [15:0] inner5_6_process_output;
  wire [15:0] inner6_6_process_output;
  wire [15:0] inner7_6_process_output;
  wire [15:0] inner8_6_process_output;
  wire [15:0] inner9_6_process_output;
  wire [15:0] inner10_6_process_output;
  wire [15:0] inner11_6_process_output;
  wire [15:0] inner12_6_process_output;
  wire [15:0] inner13_6_process_output;
  wire [15:0] inner14_6_process_output;
  wire [15:0] inner15_6_process_output;
  wire [15:0] inner0_7_process_output;
  wire [15:0] inner1_7_process_output;
  wire [15:0] inner2_7_process_output;
  wire [15:0] inner3_7_process_output;
  wire [15:0] inner4_7_process_output;
  wire [15:0] inner5_7_process_output;
  wire [15:0] inner6_7_process_output;
  wire [15:0] inner7_7_process_output;
  wire [15:0] inner8_7_process_output;
  wire [15:0] inner9_7_process_output;
  wire [15:0] inner10_7_process_output;
  wire [15:0] inner11_7_process_output;
  wire [15:0] inner12_7_process_output;
  wire [15:0] inner13_7_process_output;
  wire [15:0] inner14_7_process_output;
  wire [15:0] inner15_7_process_output;
  wire [15:0] inner0_8_process_output;
  wire [15:0] inner1_8_process_output;
  wire [15:0] inner2_8_process_output;
  wire [15:0] inner3_8_process_output;
  wire [15:0] inner4_8_process_output;
  wire [15:0] inner5_8_process_output;
  wire [15:0] inner6_8_process_output;
  wire [15:0] inner7_8_process_output;
  wire [15:0] inner8_8_process_output;
  wire [15:0] inner9_8_process_output;
  wire [15:0] inner10_8_process_output;
  wire [15:0] inner11_8_process_output;
  wire [15:0] inner12_8_process_output;
  wire [15:0] inner13_8_process_output;
  wire [15:0] inner14_8_process_output;
  wire [15:0] inner15_8_process_output;
  wire [15:0] inner0_9_process_output;
  wire [15:0] inner1_9_process_output;
  wire [15:0] inner2_9_process_output;
  wire [15:0] inner3_9_process_output;
  wire [15:0] inner4_9_process_output;
  wire [15:0] inner5_9_process_output;
  wire [15:0] inner6_9_process_output;
  wire [15:0] inner7_9_process_output;
  wire [15:0] inner8_9_process_output;
  wire [15:0] inner9_9_process_output;
  wire [15:0] inner10_9_process_output;
  wire [15:0] inner11_9_process_output;
  wire [15:0] inner12_9_process_output;
  wire [15:0] inner13_9_process_output;
  wire [15:0] inner14_9_process_output;
  wire [15:0] inner15_9_process_output;
  wire [15:0] inner0_10_process_output;
  wire [15:0] inner1_10_process_output;
  wire [15:0] inner2_10_process_output;
  wire [15:0] inner3_10_process_output;
  wire [15:0] inner4_10_process_output;
  wire [15:0] inner5_10_process_output;
  wire [15:0] inner6_10_process_output;
  wire [15:0] inner7_10_process_output;
  wire [15:0] inner8_10_process_output;
  wire [15:0] inner9_10_process_output;
  wire [15:0] inner10_10_process_output;
  wire [15:0] inner11_10_process_output;
  wire [15:0] inner12_10_process_output;
  wire [15:0] inner13_10_process_output;
  wire [15:0] inner14_10_process_output;
  wire [15:0] inner15_10_process_output;
  wire [15:0] inner0_11_process_output;
  wire [15:0] inner1_11_process_output;
  wire [15:0] inner2_11_process_output;
  wire [15:0] inner3_11_process_output;
  wire [15:0] inner4_11_process_output;
  wire [15:0] inner5_11_process_output;
  wire [15:0] inner6_11_process_output;
  wire [15:0] inner7_11_process_output;
  wire [15:0] inner8_11_process_output;
  wire [15:0] inner9_11_process_output;
  wire [15:0] inner10_11_process_output;
  wire [15:0] inner11_11_process_output;
  wire [15:0] inner12_11_process_output;
  wire [15:0] inner13_11_process_output;
  wire [15:0] inner14_11_process_output;
  wire [15:0] inner15_11_process_output;
  wire [15:0] inner0_12_process_output;
  wire [15:0] inner1_12_process_output;
  wire [15:0] inner2_12_process_output;
  wire [15:0] inner3_12_process_output;
  wire [15:0] inner4_12_process_output;
  wire [15:0] inner5_12_process_output;
  wire [15:0] inner6_12_process_output;
  wire [15:0] inner7_12_process_output;
  wire [15:0] inner8_12_process_output;
  wire [15:0] inner9_12_process_output;
  wire [15:0] inner10_12_process_output;
  wire [15:0] inner11_12_process_output;
  wire [15:0] inner12_12_process_output;
  wire [15:0] inner13_12_process_output;
  wire [15:0] inner14_12_process_output;
  wire [15:0] inner15_12_process_output;
  wire [15:0] inner0_13_process_output;
  wire [15:0] inner1_13_process_output;
  wire [15:0] inner2_13_process_output;
  wire [15:0] inner3_13_process_output;
  wire [15:0] inner4_13_process_output;
  wire [15:0] inner5_13_process_output;
  wire [15:0] inner6_13_process_output;
  wire [15:0] inner7_13_process_output;
  wire [15:0] inner8_13_process_output;
  wire [15:0] inner9_13_process_output;
  wire [15:0] inner10_13_process_output;
  wire [15:0] inner11_13_process_output;
  wire [15:0] inner12_13_process_output;
  wire [15:0] inner13_13_process_output;
  wire [15:0] inner14_13_process_output;
  wire [15:0] inner15_13_process_output;
  wire [15:0] inner0_14_process_output;
  wire [15:0] inner1_14_process_output;
  wire [15:0] inner2_14_process_output;
  wire [15:0] inner3_14_process_output;
  wire [15:0] inner4_14_process_output;
  wire [15:0] inner5_14_process_output;
  wire [15:0] inner6_14_process_output;
  wire [15:0] inner7_14_process_output;
  wire [15:0] inner8_14_process_output;
  wire [15:0] inner9_14_process_output;
  wire [15:0] inner10_14_process_output;
  wire [15:0] inner11_14_process_output;
  wire [15:0] inner12_14_process_output;
  wire [15:0] inner13_14_process_output;
  wire [15:0] inner14_14_process_output;
  wire [15:0] inner15_14_process_output;
  wire [15:0] inner0_15_process_output;
  wire [15:0] inner1_15_process_output;
  wire [15:0] inner2_15_process_output;
  wire [15:0] inner3_15_process_output;
  wire [15:0] inner4_15_process_output;
  wire [15:0] inner5_15_process_output;
  wire [15:0] inner6_15_process_output;
  wire [15:0] inner7_15_process_output;
  wire [15:0] inner8_15_process_output;
  wire [15:0] inner9_15_process_output;
  wire [15:0] inner10_15_process_output;
  wire [15:0] inner11_15_process_output;
  wire [15:0] inner12_15_process_output;
  wire [15:0] inner13_15_process_output;
  wire [15:0] inner14_15_process_output;
  wire [15:0] inner15_15_process_output;
  assign process_output = {inner15_15_process_output,inner14_15_process_output,inner13_15_process_output,inner12_15_process_output,inner11_15_process_output,inner10_15_process_output,inner9_15_process_output,inner8_15_process_output,inner7_15_process_output,inner6_15_process_output,inner5_15_process_output,inner4_15_process_output,inner3_15_process_output,inner2_15_process_output,inner1_15_process_output,inner0_15_process_output,inner15_14_process_output,inner14_14_process_output,inner13_14_process_output,inner12_14_process_output,inner11_14_process_output,inner10_14_process_output,inner9_14_process_output,inner8_14_process_output,inner7_14_process_output,inner6_14_process_output,inner5_14_process_output,inner4_14_process_output,inner3_14_process_output,inner2_14_process_output,inner1_14_process_output,inner0_14_process_output,inner15_13_process_output,inner14_13_process_output,inner13_13_process_output,inner12_13_process_output,inner11_13_process_output,inner10_13_process_output,inner9_13_process_output,inner8_13_process_output,inner7_13_process_output,inner6_13_process_output,inner5_13_process_output,inner4_13_process_output,inner3_13_process_output,inner2_13_process_output,inner1_13_process_output,inner0_13_process_output,inner15_12_process_output,inner14_12_process_output,inner13_12_process_output,inner12_12_process_output,inner11_12_process_output,inner10_12_process_output,inner9_12_process_output,inner8_12_process_output,inner7_12_process_output,inner6_12_process_output,inner5_12_process_output,inner4_12_process_output,inner3_12_process_output,inner2_12_process_output,inner1_12_process_output,inner0_12_process_output,inner15_11_process_output,inner14_11_process_output,inner13_11_process_output,inner12_11_process_output,inner11_11_process_output,inner10_11_process_output,inner9_11_process_output,inner8_11_process_output,inner7_11_process_output,inner6_11_process_output,inner5_11_process_output,inner4_11_process_output,inner3_11_process_output,inner2_11_process_output,inner1_11_process_output,inner0_11_process_output,inner15_10_process_output,inner14_10_process_output,inner13_10_process_output,inner12_10_process_output,inner11_10_process_output,inner10_10_process_output,inner9_10_process_output,inner8_10_process_output,inner7_10_process_output,inner6_10_process_output,inner5_10_process_output,inner4_10_process_output,inner3_10_process_output,inner2_10_process_output,inner1_10_process_output,inner0_10_process_output,inner15_9_process_output,inner14_9_process_output,inner13_9_process_output,inner12_9_process_output,inner11_9_process_output,inner10_9_process_output,inner9_9_process_output,inner8_9_process_output,inner7_9_process_output,inner6_9_process_output,inner5_9_process_output,inner4_9_process_output,inner3_9_process_output,inner2_9_process_output,inner1_9_process_output,inner0_9_process_output,inner15_8_process_output,inner14_8_process_output,inner13_8_process_output,inner12_8_process_output,inner11_8_process_output,inner10_8_process_output,inner9_8_process_output,inner8_8_process_output,inner7_8_process_output,inner6_8_process_output,inner5_8_process_output,inner4_8_process_output,inner3_8_process_output,inner2_8_process_output,inner1_8_process_output,inner0_8_process_output,inner15_7_process_output,inner14_7_process_output,inner13_7_process_output,inner12_7_process_output,inner11_7_process_output,inner10_7_process_output,inner9_7_process_output,inner8_7_process_output,inner7_7_process_output,inner6_7_process_output,inner5_7_process_output,inner4_7_process_output,inner3_7_process_output,inner2_7_process_output,inner1_7_process_output,inner0_7_process_output,inner15_6_process_output,inner14_6_process_output,inner13_6_process_output,inner12_6_process_output,inner11_6_process_output,inner10_6_process_output,inner9_6_process_output,inner8_6_process_output,inner7_6_process_output,inner6_6_process_output,inner5_6_process_output,inner4_6_process_output,inner3_6_process_output,inner2_6_process_output,inner1_6_process_output,inner0_6_process_output,inner15_5_process_output,inner14_5_process_output,inner13_5_process_output,inner12_5_process_output,inner11_5_process_output,inner10_5_process_output,inner9_5_process_output,inner8_5_process_output,inner7_5_process_output,inner6_5_process_output,inner5_5_process_output,inner4_5_process_output,inner3_5_process_output,inner2_5_process_output,inner1_5_process_output,inner0_5_process_output,inner15_4_process_output,inner14_4_process_output,inner13_4_process_output,inner12_4_process_output,inner11_4_process_output,inner10_4_process_output,inner9_4_process_output,inner8_4_process_output,inner7_4_process_output,inner6_4_process_output,inner5_4_process_output,inner4_4_process_output,inner3_4_process_output,inner2_4_process_output,inner1_4_process_output,inner0_4_process_output,inner15_3_process_output,inner14_3_process_output,inner13_3_process_output,inner12_3_process_output,inner11_3_process_output,inner10_3_process_output,inner9_3_process_output,inner8_3_process_output,inner7_3_process_output,inner6_3_process_output,inner5_3_process_output,inner4_3_process_output,inner3_3_process_output,inner2_3_process_output,inner1_3_process_output,inner0_3_process_output,inner15_2_process_output,inner14_2_process_output,inner13_2_process_output,inner12_2_process_output,inner11_2_process_output,inner10_2_process_output,inner9_2_process_output,inner8_2_process_output,inner7_2_process_output,inner6_2_process_output,inner5_2_process_output,inner4_2_process_output,inner3_2_process_output,inner2_2_process_output,inner1_2_process_output,inner0_2_process_output,inner15_1_process_output,inner14_1_process_output,inner13_1_process_output,inner12_1_process_output,inner11_1_process_output,inner10_1_process_output,inner9_1_process_output,inner8_1_process_output,inner7_1_process_output,inner6_1_process_output,inner5_1_process_output,inner4_1_process_output,inner3_1_process_output,inner2_1_process_output,inner1_1_process_output,inner0_1_process_output,inner15_0_process_output,inner14_0_process_output,inner13_0_process_output,inner12_0_process_output,inner11_0_process_output,inner10_0_process_output,inner9_0_process_output,inner8_0_process_output,inner7_0_process_output,inner6_0_process_output,inner5_0_process_output,inner4_0_process_output,inner3_0_process_output,inner2_0_process_output,inner1_0_process_output,inner0_0_process_output};
  // function: process pure=true delay=3
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner0_0"})) inner0_0(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[15:0]})), .process_output(inner0_0_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner1_0"})) inner1_0(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[31:16]})), .process_output(inner1_0_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner2_0"})) inner2_0(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[47:32]})), .process_output(inner2_0_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner3_0"})) inner3_0(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[63:48]})), .process_output(inner3_0_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner4_0"})) inner4_0(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[79:64]})), .process_output(inner4_0_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner5_0"})) inner5_0(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[95:80]})), .process_output(inner5_0_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner6_0"})) inner6_0(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[111:96]})), .process_output(inner6_0_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner7_0"})) inner7_0(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[127:112]})), .process_output(inner7_0_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner8_0"})) inner8_0(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[143:128]})), .process_output(inner8_0_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner9_0"})) inner9_0(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[159:144]})), .process_output(inner9_0_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner10_0"})) inner10_0(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[175:160]})), .process_output(inner10_0_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner11_0"})) inner11_0(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[191:176]})), .process_output(inner11_0_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner12_0"})) inner12_0(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[207:192]})), .process_output(inner12_0_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner13_0"})) inner13_0(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[223:208]})), .process_output(inner13_0_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner14_0"})) inner14_0(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[239:224]})), .process_output(inner14_0_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner15_0"})) inner15_0(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[255:240]})), .process_output(inner15_0_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner0_1"})) inner0_1(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[271:256]})), .process_output(inner0_1_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner1_1"})) inner1_1(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[287:272]})), .process_output(inner1_1_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner2_1"})) inner2_1(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[303:288]})), .process_output(inner2_1_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner3_1"})) inner3_1(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[319:304]})), .process_output(inner3_1_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner4_1"})) inner4_1(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[335:320]})), .process_output(inner4_1_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner5_1"})) inner5_1(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[351:336]})), .process_output(inner5_1_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner6_1"})) inner6_1(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[367:352]})), .process_output(inner6_1_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner7_1"})) inner7_1(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[383:368]})), .process_output(inner7_1_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner8_1"})) inner8_1(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[399:384]})), .process_output(inner8_1_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner9_1"})) inner9_1(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[415:400]})), .process_output(inner9_1_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner10_1"})) inner10_1(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[431:416]})), .process_output(inner10_1_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner11_1"})) inner11_1(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[447:432]})), .process_output(inner11_1_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner12_1"})) inner12_1(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[463:448]})), .process_output(inner12_1_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner13_1"})) inner13_1(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[479:464]})), .process_output(inner13_1_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner14_1"})) inner14_1(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[495:480]})), .process_output(inner14_1_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner15_1"})) inner15_1(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[511:496]})), .process_output(inner15_1_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner0_2"})) inner0_2(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[527:512]})), .process_output(inner0_2_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner1_2"})) inner1_2(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[543:528]})), .process_output(inner1_2_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner2_2"})) inner2_2(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[559:544]})), .process_output(inner2_2_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner3_2"})) inner3_2(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[575:560]})), .process_output(inner3_2_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner4_2"})) inner4_2(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[591:576]})), .process_output(inner4_2_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner5_2"})) inner5_2(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[607:592]})), .process_output(inner5_2_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner6_2"})) inner6_2(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[623:608]})), .process_output(inner6_2_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner7_2"})) inner7_2(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[639:624]})), .process_output(inner7_2_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner8_2"})) inner8_2(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[655:640]})), .process_output(inner8_2_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner9_2"})) inner9_2(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[671:656]})), .process_output(inner9_2_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner10_2"})) inner10_2(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[687:672]})), .process_output(inner10_2_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner11_2"})) inner11_2(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[703:688]})), .process_output(inner11_2_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner12_2"})) inner12_2(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[719:704]})), .process_output(inner12_2_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner13_2"})) inner13_2(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[735:720]})), .process_output(inner13_2_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner14_2"})) inner14_2(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[751:736]})), .process_output(inner14_2_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner15_2"})) inner15_2(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[767:752]})), .process_output(inner15_2_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner0_3"})) inner0_3(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[783:768]})), .process_output(inner0_3_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner1_3"})) inner1_3(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[799:784]})), .process_output(inner1_3_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner2_3"})) inner2_3(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[815:800]})), .process_output(inner2_3_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner3_3"})) inner3_3(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[831:816]})), .process_output(inner3_3_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner4_3"})) inner4_3(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[847:832]})), .process_output(inner4_3_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner5_3"})) inner5_3(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[863:848]})), .process_output(inner5_3_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner6_3"})) inner6_3(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[879:864]})), .process_output(inner6_3_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner7_3"})) inner7_3(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[895:880]})), .process_output(inner7_3_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner8_3"})) inner8_3(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[911:896]})), .process_output(inner8_3_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner9_3"})) inner9_3(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[927:912]})), .process_output(inner9_3_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner10_3"})) inner10_3(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[943:928]})), .process_output(inner10_3_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner11_3"})) inner11_3(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[959:944]})), .process_output(inner11_3_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner12_3"})) inner12_3(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[975:960]})), .process_output(inner12_3_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner13_3"})) inner13_3(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[991:976]})), .process_output(inner13_3_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner14_3"})) inner14_3(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1007:992]})), .process_output(inner14_3_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner15_3"})) inner15_3(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1023:1008]})), .process_output(inner15_3_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner0_4"})) inner0_4(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1039:1024]})), .process_output(inner0_4_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner1_4"})) inner1_4(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1055:1040]})), .process_output(inner1_4_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner2_4"})) inner2_4(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1071:1056]})), .process_output(inner2_4_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner3_4"})) inner3_4(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1087:1072]})), .process_output(inner3_4_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner4_4"})) inner4_4(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1103:1088]})), .process_output(inner4_4_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner5_4"})) inner5_4(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1119:1104]})), .process_output(inner5_4_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner6_4"})) inner6_4(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1135:1120]})), .process_output(inner6_4_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner7_4"})) inner7_4(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1151:1136]})), .process_output(inner7_4_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner8_4"})) inner8_4(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1167:1152]})), .process_output(inner8_4_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner9_4"})) inner9_4(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1183:1168]})), .process_output(inner9_4_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner10_4"})) inner10_4(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1199:1184]})), .process_output(inner10_4_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner11_4"})) inner11_4(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1215:1200]})), .process_output(inner11_4_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner12_4"})) inner12_4(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1231:1216]})), .process_output(inner12_4_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner13_4"})) inner13_4(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1247:1232]})), .process_output(inner13_4_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner14_4"})) inner14_4(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1263:1248]})), .process_output(inner14_4_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner15_4"})) inner15_4(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1279:1264]})), .process_output(inner15_4_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner0_5"})) inner0_5(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1295:1280]})), .process_output(inner0_5_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner1_5"})) inner1_5(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1311:1296]})), .process_output(inner1_5_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner2_5"})) inner2_5(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1327:1312]})), .process_output(inner2_5_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner3_5"})) inner3_5(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1343:1328]})), .process_output(inner3_5_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner4_5"})) inner4_5(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1359:1344]})), .process_output(inner4_5_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner5_5"})) inner5_5(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1375:1360]})), .process_output(inner5_5_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner6_5"})) inner6_5(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1391:1376]})), .process_output(inner6_5_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner7_5"})) inner7_5(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1407:1392]})), .process_output(inner7_5_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner8_5"})) inner8_5(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1423:1408]})), .process_output(inner8_5_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner9_5"})) inner9_5(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1439:1424]})), .process_output(inner9_5_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner10_5"})) inner10_5(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1455:1440]})), .process_output(inner10_5_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner11_5"})) inner11_5(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1471:1456]})), .process_output(inner11_5_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner12_5"})) inner12_5(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1487:1472]})), .process_output(inner12_5_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner13_5"})) inner13_5(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1503:1488]})), .process_output(inner13_5_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner14_5"})) inner14_5(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1519:1504]})), .process_output(inner14_5_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner15_5"})) inner15_5(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1535:1520]})), .process_output(inner15_5_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner0_6"})) inner0_6(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1551:1536]})), .process_output(inner0_6_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner1_6"})) inner1_6(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1567:1552]})), .process_output(inner1_6_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner2_6"})) inner2_6(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1583:1568]})), .process_output(inner2_6_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner3_6"})) inner3_6(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1599:1584]})), .process_output(inner3_6_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner4_6"})) inner4_6(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1615:1600]})), .process_output(inner4_6_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner5_6"})) inner5_6(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1631:1616]})), .process_output(inner5_6_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner6_6"})) inner6_6(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1647:1632]})), .process_output(inner6_6_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner7_6"})) inner7_6(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1663:1648]})), .process_output(inner7_6_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner8_6"})) inner8_6(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1679:1664]})), .process_output(inner8_6_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner9_6"})) inner9_6(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1695:1680]})), .process_output(inner9_6_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner10_6"})) inner10_6(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1711:1696]})), .process_output(inner10_6_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner11_6"})) inner11_6(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1727:1712]})), .process_output(inner11_6_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner12_6"})) inner12_6(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1743:1728]})), .process_output(inner12_6_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner13_6"})) inner13_6(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1759:1744]})), .process_output(inner13_6_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner14_6"})) inner14_6(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1775:1760]})), .process_output(inner14_6_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner15_6"})) inner15_6(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1791:1776]})), .process_output(inner15_6_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner0_7"})) inner0_7(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1807:1792]})), .process_output(inner0_7_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner1_7"})) inner1_7(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1823:1808]})), .process_output(inner1_7_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner2_7"})) inner2_7(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1839:1824]})), .process_output(inner2_7_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner3_7"})) inner3_7(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1855:1840]})), .process_output(inner3_7_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner4_7"})) inner4_7(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1871:1856]})), .process_output(inner4_7_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner5_7"})) inner5_7(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1887:1872]})), .process_output(inner5_7_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner6_7"})) inner6_7(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1903:1888]})), .process_output(inner6_7_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner7_7"})) inner7_7(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1919:1904]})), .process_output(inner7_7_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner8_7"})) inner8_7(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1935:1920]})), .process_output(inner8_7_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner9_7"})) inner9_7(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1951:1936]})), .process_output(inner9_7_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner10_7"})) inner10_7(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1967:1952]})), .process_output(inner10_7_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner11_7"})) inner11_7(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1983:1968]})), .process_output(inner11_7_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner12_7"})) inner12_7(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[1999:1984]})), .process_output(inner12_7_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner13_7"})) inner13_7(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2015:2000]})), .process_output(inner13_7_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner14_7"})) inner14_7(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2031:2016]})), .process_output(inner14_7_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner15_7"})) inner15_7(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2047:2032]})), .process_output(inner15_7_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner0_8"})) inner0_8(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2063:2048]})), .process_output(inner0_8_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner1_8"})) inner1_8(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2079:2064]})), .process_output(inner1_8_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner2_8"})) inner2_8(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2095:2080]})), .process_output(inner2_8_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner3_8"})) inner3_8(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2111:2096]})), .process_output(inner3_8_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner4_8"})) inner4_8(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2127:2112]})), .process_output(inner4_8_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner5_8"})) inner5_8(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2143:2128]})), .process_output(inner5_8_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner6_8"})) inner6_8(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2159:2144]})), .process_output(inner6_8_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner7_8"})) inner7_8(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2175:2160]})), .process_output(inner7_8_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner8_8"})) inner8_8(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2191:2176]})), .process_output(inner8_8_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner9_8"})) inner9_8(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2207:2192]})), .process_output(inner9_8_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner10_8"})) inner10_8(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2223:2208]})), .process_output(inner10_8_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner11_8"})) inner11_8(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2239:2224]})), .process_output(inner11_8_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner12_8"})) inner12_8(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2255:2240]})), .process_output(inner12_8_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner13_8"})) inner13_8(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2271:2256]})), .process_output(inner13_8_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner14_8"})) inner14_8(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2287:2272]})), .process_output(inner14_8_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner15_8"})) inner15_8(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2303:2288]})), .process_output(inner15_8_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner0_9"})) inner0_9(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2319:2304]})), .process_output(inner0_9_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner1_9"})) inner1_9(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2335:2320]})), .process_output(inner1_9_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner2_9"})) inner2_9(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2351:2336]})), .process_output(inner2_9_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner3_9"})) inner3_9(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2367:2352]})), .process_output(inner3_9_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner4_9"})) inner4_9(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2383:2368]})), .process_output(inner4_9_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner5_9"})) inner5_9(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2399:2384]})), .process_output(inner5_9_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner6_9"})) inner6_9(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2415:2400]})), .process_output(inner6_9_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner7_9"})) inner7_9(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2431:2416]})), .process_output(inner7_9_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner8_9"})) inner8_9(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2447:2432]})), .process_output(inner8_9_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner9_9"})) inner9_9(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2463:2448]})), .process_output(inner9_9_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner10_9"})) inner10_9(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2479:2464]})), .process_output(inner10_9_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner11_9"})) inner11_9(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2495:2480]})), .process_output(inner11_9_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner12_9"})) inner12_9(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2511:2496]})), .process_output(inner12_9_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner13_9"})) inner13_9(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2527:2512]})), .process_output(inner13_9_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner14_9"})) inner14_9(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2543:2528]})), .process_output(inner14_9_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner15_9"})) inner15_9(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2559:2544]})), .process_output(inner15_9_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner0_10"})) inner0_10(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2575:2560]})), .process_output(inner0_10_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner1_10"})) inner1_10(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2591:2576]})), .process_output(inner1_10_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner2_10"})) inner2_10(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2607:2592]})), .process_output(inner2_10_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner3_10"})) inner3_10(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2623:2608]})), .process_output(inner3_10_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner4_10"})) inner4_10(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2639:2624]})), .process_output(inner4_10_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner5_10"})) inner5_10(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2655:2640]})), .process_output(inner5_10_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner6_10"})) inner6_10(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2671:2656]})), .process_output(inner6_10_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner7_10"})) inner7_10(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2687:2672]})), .process_output(inner7_10_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner8_10"})) inner8_10(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2703:2688]})), .process_output(inner8_10_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner9_10"})) inner9_10(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2719:2704]})), .process_output(inner9_10_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner10_10"})) inner10_10(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2735:2720]})), .process_output(inner10_10_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner11_10"})) inner11_10(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2751:2736]})), .process_output(inner11_10_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner12_10"})) inner12_10(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2767:2752]})), .process_output(inner12_10_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner13_10"})) inner13_10(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2783:2768]})), .process_output(inner13_10_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner14_10"})) inner14_10(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2799:2784]})), .process_output(inner14_10_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner15_10"})) inner15_10(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2815:2800]})), .process_output(inner15_10_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner0_11"})) inner0_11(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2831:2816]})), .process_output(inner0_11_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner1_11"})) inner1_11(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2847:2832]})), .process_output(inner1_11_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner2_11"})) inner2_11(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2863:2848]})), .process_output(inner2_11_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner3_11"})) inner3_11(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2879:2864]})), .process_output(inner3_11_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner4_11"})) inner4_11(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2895:2880]})), .process_output(inner4_11_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner5_11"})) inner5_11(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2911:2896]})), .process_output(inner5_11_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner6_11"})) inner6_11(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2927:2912]})), .process_output(inner6_11_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner7_11"})) inner7_11(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2943:2928]})), .process_output(inner7_11_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner8_11"})) inner8_11(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2959:2944]})), .process_output(inner8_11_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner9_11"})) inner9_11(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2975:2960]})), .process_output(inner9_11_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner10_11"})) inner10_11(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[2991:2976]})), .process_output(inner10_11_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner11_11"})) inner11_11(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3007:2992]})), .process_output(inner11_11_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner12_11"})) inner12_11(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3023:3008]})), .process_output(inner12_11_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner13_11"})) inner13_11(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3039:3024]})), .process_output(inner13_11_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner14_11"})) inner14_11(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3055:3040]})), .process_output(inner14_11_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner15_11"})) inner15_11(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3071:3056]})), .process_output(inner15_11_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner0_12"})) inner0_12(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3087:3072]})), .process_output(inner0_12_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner1_12"})) inner1_12(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3103:3088]})), .process_output(inner1_12_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner2_12"})) inner2_12(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3119:3104]})), .process_output(inner2_12_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner3_12"})) inner3_12(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3135:3120]})), .process_output(inner3_12_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner4_12"})) inner4_12(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3151:3136]})), .process_output(inner4_12_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner5_12"})) inner5_12(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3167:3152]})), .process_output(inner5_12_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner6_12"})) inner6_12(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3183:3168]})), .process_output(inner6_12_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner7_12"})) inner7_12(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3199:3184]})), .process_output(inner7_12_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner8_12"})) inner8_12(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3215:3200]})), .process_output(inner8_12_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner9_12"})) inner9_12(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3231:3216]})), .process_output(inner9_12_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner10_12"})) inner10_12(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3247:3232]})), .process_output(inner10_12_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner11_12"})) inner11_12(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3263:3248]})), .process_output(inner11_12_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner12_12"})) inner12_12(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3279:3264]})), .process_output(inner12_12_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner13_12"})) inner13_12(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3295:3280]})), .process_output(inner13_12_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner14_12"})) inner14_12(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3311:3296]})), .process_output(inner14_12_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner15_12"})) inner15_12(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3327:3312]})), .process_output(inner15_12_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner0_13"})) inner0_13(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3343:3328]})), .process_output(inner0_13_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner1_13"})) inner1_13(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3359:3344]})), .process_output(inner1_13_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner2_13"})) inner2_13(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3375:3360]})), .process_output(inner2_13_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner3_13"})) inner3_13(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3391:3376]})), .process_output(inner3_13_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner4_13"})) inner4_13(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3407:3392]})), .process_output(inner4_13_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner5_13"})) inner5_13(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3423:3408]})), .process_output(inner5_13_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner6_13"})) inner6_13(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3439:3424]})), .process_output(inner6_13_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner7_13"})) inner7_13(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3455:3440]})), .process_output(inner7_13_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner8_13"})) inner8_13(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3471:3456]})), .process_output(inner8_13_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner9_13"})) inner9_13(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3487:3472]})), .process_output(inner9_13_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner10_13"})) inner10_13(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3503:3488]})), .process_output(inner10_13_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner11_13"})) inner11_13(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3519:3504]})), .process_output(inner11_13_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner12_13"})) inner12_13(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3535:3520]})), .process_output(inner12_13_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner13_13"})) inner13_13(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3551:3536]})), .process_output(inner13_13_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner14_13"})) inner14_13(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3567:3552]})), .process_output(inner14_13_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner15_13"})) inner15_13(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3583:3568]})), .process_output(inner15_13_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner0_14"})) inner0_14(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3599:3584]})), .process_output(inner0_14_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner1_14"})) inner1_14(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3615:3600]})), .process_output(inner1_14_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner2_14"})) inner2_14(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3631:3616]})), .process_output(inner2_14_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner3_14"})) inner3_14(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3647:3632]})), .process_output(inner3_14_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner4_14"})) inner4_14(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3663:3648]})), .process_output(inner4_14_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner5_14"})) inner5_14(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3679:3664]})), .process_output(inner5_14_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner6_14"})) inner6_14(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3695:3680]})), .process_output(inner6_14_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner7_14"})) inner7_14(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3711:3696]})), .process_output(inner7_14_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner8_14"})) inner8_14(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3727:3712]})), .process_output(inner8_14_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner9_14"})) inner9_14(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3743:3728]})), .process_output(inner9_14_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner10_14"})) inner10_14(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3759:3744]})), .process_output(inner10_14_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner11_14"})) inner11_14(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3775:3760]})), .process_output(inner11_14_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner12_14"})) inner12_14(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3791:3776]})), .process_output(inner12_14_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner13_14"})) inner13_14(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3807:3792]})), .process_output(inner13_14_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner14_14"})) inner14_14(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3823:3808]})), .process_output(inner14_14_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner15_14"})) inner15_14(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3839:3824]})), .process_output(inner15_14_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner0_15"})) inner0_15(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3855:3840]})), .process_output(inner0_15_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner1_15"})) inner1_15(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3871:3856]})), .process_output(inner1_15_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner2_15"})) inner2_15(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3887:3872]})), .process_output(inner2_15_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner3_15"})) inner3_15(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3903:3888]})), .process_output(inner3_15_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner4_15"})) inner4_15(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3919:3904]})), .process_output(inner4_15_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner5_15"})) inner5_15(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3935:3920]})), .process_output(inner5_15_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner6_15"})) inner6_15(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3951:3936]})), .process_output(inner6_15_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner7_15"})) inner7_15(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3967:3952]})), .process_output(inner7_15_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner8_15"})) inner8_15(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3983:3968]})), .process_output(inner8_15_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner9_15"})) inner9_15(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[3999:3984]})), .process_output(inner9_15_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner10_15"})) inner10_15(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[4015:4000]})), .process_output(inner10_15_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner11_15"})) inner11_15(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[4031:4016]})), .process_output(inner11_15_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner12_15"})) inner12_15(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[4047:4032]})), .process_output(inner12_15_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner13_15"})) inner13_15(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[4063:4048]})), .process_output(inner13_15_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner14_15"})) inner14_15(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[4079:4064]})), .process_output(inner14_15_process_output));
  absoluteDiff #(.INSTANCE_NAME({INSTANCE_NAME,"_inner15_15"})) inner15_15(.CLK(CLK), .process_CE(process_CE), .abs_inp(({process_input[4095:4080]})), .process_output(inner15_15_process_output));
endmodule

module ABS_SUM(input CLK, input process_CE, input [31:0] sum_inp, output [15:0] process_output);
parameter INSTANCE_NAME="INST";
  reg [16:0] unnamedbinop30140_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop30140_delay1_validunnamednull0_CEprocess_CE <= {({1'b0,(sum_inp[15:0])}+{1'b0,(sum_inp[31:16])})}; end end
  assign process_output = {unnamedbinop30140_delay1_validunnamednull0_CEprocess_CE[15:0]};
  // function: process pure=true delay=1
endmodule

module reduce_ABS_SUM_W16_H16(input CLK, input process_CE, input [4095:0] process_input, output [15:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] inner0_process_output;
  wire [15:0] inner1_process_output;
  wire [15:0] inner128_process_output;
  wire [15:0] inner2_process_output;
  wire [15:0] inner3_process_output;
  wire [15:0] inner129_process_output;
  wire [15:0] inner192_process_output;
  wire [15:0] inner4_process_output;
  wire [15:0] inner5_process_output;
  wire [15:0] inner130_process_output;
  wire [15:0] inner6_process_output;
  wire [15:0] inner7_process_output;
  wire [15:0] inner131_process_output;
  wire [15:0] inner193_process_output;
  wire [15:0] inner224_process_output;
  wire [15:0] inner8_process_output;
  wire [15:0] inner9_process_output;
  wire [15:0] inner132_process_output;
  wire [15:0] inner10_process_output;
  wire [15:0] inner11_process_output;
  wire [15:0] inner133_process_output;
  wire [15:0] inner194_process_output;
  wire [15:0] inner12_process_output;
  wire [15:0] inner13_process_output;
  wire [15:0] inner134_process_output;
  wire [15:0] inner14_process_output;
  wire [15:0] inner15_process_output;
  wire [15:0] inner135_process_output;
  wire [15:0] inner195_process_output;
  wire [15:0] inner225_process_output;
  wire [15:0] inner240_process_output;
  wire [15:0] inner16_process_output;
  wire [15:0] inner17_process_output;
  wire [15:0] inner136_process_output;
  wire [15:0] inner18_process_output;
  wire [15:0] inner19_process_output;
  wire [15:0] inner137_process_output;
  wire [15:0] inner196_process_output;
  wire [15:0] inner20_process_output;
  wire [15:0] inner21_process_output;
  wire [15:0] inner138_process_output;
  wire [15:0] inner22_process_output;
  wire [15:0] inner23_process_output;
  wire [15:0] inner139_process_output;
  wire [15:0] inner197_process_output;
  wire [15:0] inner226_process_output;
  wire [15:0] inner24_process_output;
  wire [15:0] inner25_process_output;
  wire [15:0] inner140_process_output;
  wire [15:0] inner26_process_output;
  wire [15:0] inner27_process_output;
  wire [15:0] inner141_process_output;
  wire [15:0] inner198_process_output;
  wire [15:0] inner28_process_output;
  wire [15:0] inner29_process_output;
  wire [15:0] inner142_process_output;
  wire [15:0] inner30_process_output;
  wire [15:0] inner31_process_output;
  wire [15:0] inner143_process_output;
  wire [15:0] inner199_process_output;
  wire [15:0] inner227_process_output;
  wire [15:0] inner241_process_output;
  wire [15:0] inner248_process_output;
  wire [15:0] inner32_process_output;
  wire [15:0] inner33_process_output;
  wire [15:0] inner144_process_output;
  wire [15:0] inner34_process_output;
  wire [15:0] inner35_process_output;
  wire [15:0] inner145_process_output;
  wire [15:0] inner200_process_output;
  wire [15:0] inner36_process_output;
  wire [15:0] inner37_process_output;
  wire [15:0] inner146_process_output;
  wire [15:0] inner38_process_output;
  wire [15:0] inner39_process_output;
  wire [15:0] inner147_process_output;
  wire [15:0] inner201_process_output;
  wire [15:0] inner228_process_output;
  wire [15:0] inner40_process_output;
  wire [15:0] inner41_process_output;
  wire [15:0] inner148_process_output;
  wire [15:0] inner42_process_output;
  wire [15:0] inner43_process_output;
  wire [15:0] inner149_process_output;
  wire [15:0] inner202_process_output;
  wire [15:0] inner44_process_output;
  wire [15:0] inner45_process_output;
  wire [15:0] inner150_process_output;
  wire [15:0] inner46_process_output;
  wire [15:0] inner47_process_output;
  wire [15:0] inner151_process_output;
  wire [15:0] inner203_process_output;
  wire [15:0] inner229_process_output;
  wire [15:0] inner242_process_output;
  wire [15:0] inner48_process_output;
  wire [15:0] inner49_process_output;
  wire [15:0] inner152_process_output;
  wire [15:0] inner50_process_output;
  wire [15:0] inner51_process_output;
  wire [15:0] inner153_process_output;
  wire [15:0] inner204_process_output;
  wire [15:0] inner52_process_output;
  wire [15:0] inner53_process_output;
  wire [15:0] inner154_process_output;
  wire [15:0] inner54_process_output;
  wire [15:0] inner55_process_output;
  wire [15:0] inner155_process_output;
  wire [15:0] inner205_process_output;
  wire [15:0] inner230_process_output;
  wire [15:0] inner56_process_output;
  wire [15:0] inner57_process_output;
  wire [15:0] inner156_process_output;
  wire [15:0] inner58_process_output;
  wire [15:0] inner59_process_output;
  wire [15:0] inner157_process_output;
  wire [15:0] inner206_process_output;
  wire [15:0] inner60_process_output;
  wire [15:0] inner61_process_output;
  wire [15:0] inner158_process_output;
  wire [15:0] inner62_process_output;
  wire [15:0] inner63_process_output;
  wire [15:0] inner159_process_output;
  wire [15:0] inner207_process_output;
  wire [15:0] inner231_process_output;
  wire [15:0] inner243_process_output;
  wire [15:0] inner249_process_output;
  wire [15:0] inner252_process_output;
  wire [15:0] inner64_process_output;
  wire [15:0] inner65_process_output;
  wire [15:0] inner160_process_output;
  wire [15:0] inner66_process_output;
  wire [15:0] inner67_process_output;
  wire [15:0] inner161_process_output;
  wire [15:0] inner208_process_output;
  wire [15:0] inner68_process_output;
  wire [15:0] inner69_process_output;
  wire [15:0] inner162_process_output;
  wire [15:0] inner70_process_output;
  wire [15:0] inner71_process_output;
  wire [15:0] inner163_process_output;
  wire [15:0] inner209_process_output;
  wire [15:0] inner232_process_output;
  wire [15:0] inner72_process_output;
  wire [15:0] inner73_process_output;
  wire [15:0] inner164_process_output;
  wire [15:0] inner74_process_output;
  wire [15:0] inner75_process_output;
  wire [15:0] inner165_process_output;
  wire [15:0] inner210_process_output;
  wire [15:0] inner76_process_output;
  wire [15:0] inner77_process_output;
  wire [15:0] inner166_process_output;
  wire [15:0] inner78_process_output;
  wire [15:0] inner79_process_output;
  wire [15:0] inner167_process_output;
  wire [15:0] inner211_process_output;
  wire [15:0] inner233_process_output;
  wire [15:0] inner244_process_output;
  wire [15:0] inner80_process_output;
  wire [15:0] inner81_process_output;
  wire [15:0] inner168_process_output;
  wire [15:0] inner82_process_output;
  wire [15:0] inner83_process_output;
  wire [15:0] inner169_process_output;
  wire [15:0] inner212_process_output;
  wire [15:0] inner84_process_output;
  wire [15:0] inner85_process_output;
  wire [15:0] inner170_process_output;
  wire [15:0] inner86_process_output;
  wire [15:0] inner87_process_output;
  wire [15:0] inner171_process_output;
  wire [15:0] inner213_process_output;
  wire [15:0] inner234_process_output;
  wire [15:0] inner88_process_output;
  wire [15:0] inner89_process_output;
  wire [15:0] inner172_process_output;
  wire [15:0] inner90_process_output;
  wire [15:0] inner91_process_output;
  wire [15:0] inner173_process_output;
  wire [15:0] inner214_process_output;
  wire [15:0] inner92_process_output;
  wire [15:0] inner93_process_output;
  wire [15:0] inner174_process_output;
  wire [15:0] inner94_process_output;
  wire [15:0] inner95_process_output;
  wire [15:0] inner175_process_output;
  wire [15:0] inner215_process_output;
  wire [15:0] inner235_process_output;
  wire [15:0] inner245_process_output;
  wire [15:0] inner250_process_output;
  wire [15:0] inner96_process_output;
  wire [15:0] inner97_process_output;
  wire [15:0] inner176_process_output;
  wire [15:0] inner98_process_output;
  wire [15:0] inner99_process_output;
  wire [15:0] inner177_process_output;
  wire [15:0] inner216_process_output;
  wire [15:0] inner100_process_output;
  wire [15:0] inner101_process_output;
  wire [15:0] inner178_process_output;
  wire [15:0] inner102_process_output;
  wire [15:0] inner103_process_output;
  wire [15:0] inner179_process_output;
  wire [15:0] inner217_process_output;
  wire [15:0] inner236_process_output;
  wire [15:0] inner104_process_output;
  wire [15:0] inner105_process_output;
  wire [15:0] inner180_process_output;
  wire [15:0] inner106_process_output;
  wire [15:0] inner107_process_output;
  wire [15:0] inner181_process_output;
  wire [15:0] inner218_process_output;
  wire [15:0] inner108_process_output;
  wire [15:0] inner109_process_output;
  wire [15:0] inner182_process_output;
  wire [15:0] inner110_process_output;
  wire [15:0] inner111_process_output;
  wire [15:0] inner183_process_output;
  wire [15:0] inner219_process_output;
  wire [15:0] inner237_process_output;
  wire [15:0] inner246_process_output;
  wire [15:0] inner112_process_output;
  wire [15:0] inner113_process_output;
  wire [15:0] inner184_process_output;
  wire [15:0] inner114_process_output;
  wire [15:0] inner115_process_output;
  wire [15:0] inner185_process_output;
  wire [15:0] inner220_process_output;
  wire [15:0] inner116_process_output;
  wire [15:0] inner117_process_output;
  wire [15:0] inner186_process_output;
  wire [15:0] inner118_process_output;
  wire [15:0] inner119_process_output;
  wire [15:0] inner187_process_output;
  wire [15:0] inner221_process_output;
  wire [15:0] inner238_process_output;
  wire [15:0] inner120_process_output;
  wire [15:0] inner121_process_output;
  wire [15:0] inner188_process_output;
  wire [15:0] inner122_process_output;
  wire [15:0] inner123_process_output;
  wire [15:0] inner189_process_output;
  wire [15:0] inner222_process_output;
  wire [15:0] inner124_process_output;
  wire [15:0] inner125_process_output;
  wire [15:0] inner190_process_output;
  wire [15:0] inner126_process_output;
  wire [15:0] inner127_process_output;
  wire [15:0] inner191_process_output;
  wire [15:0] inner223_process_output;
  wire [15:0] inner239_process_output;
  wire [15:0] inner247_process_output;
  wire [15:0] inner251_process_output;
  wire [15:0] inner253_process_output;
  wire [15:0] inner254_process_output;
  assign process_output = inner254_process_output;
  // function: process pure=true delay=8
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner0"})) inner0(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[31:16]}),({process_input[15:0]})}), .process_output(inner0_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner1"})) inner1(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[63:48]}),({process_input[47:32]})}), .process_output(inner1_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner2"})) inner2(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[95:80]}),({process_input[79:64]})}), .process_output(inner2_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner3"})) inner3(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[127:112]}),({process_input[111:96]})}), .process_output(inner3_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner4"})) inner4(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[159:144]}),({process_input[143:128]})}), .process_output(inner4_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner5"})) inner5(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[191:176]}),({process_input[175:160]})}), .process_output(inner5_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner6"})) inner6(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[223:208]}),({process_input[207:192]})}), .process_output(inner6_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner7"})) inner7(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[255:240]}),({process_input[239:224]})}), .process_output(inner7_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner8"})) inner8(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[287:272]}),({process_input[271:256]})}), .process_output(inner8_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner9"})) inner9(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[319:304]}),({process_input[303:288]})}), .process_output(inner9_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner10"})) inner10(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[351:336]}),({process_input[335:320]})}), .process_output(inner10_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner11"})) inner11(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[383:368]}),({process_input[367:352]})}), .process_output(inner11_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner12"})) inner12(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[415:400]}),({process_input[399:384]})}), .process_output(inner12_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner13"})) inner13(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[447:432]}),({process_input[431:416]})}), .process_output(inner13_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner14"})) inner14(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[479:464]}),({process_input[463:448]})}), .process_output(inner14_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner15"})) inner15(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[511:496]}),({process_input[495:480]})}), .process_output(inner15_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner16"})) inner16(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[543:528]}),({process_input[527:512]})}), .process_output(inner16_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner17"})) inner17(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[575:560]}),({process_input[559:544]})}), .process_output(inner17_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner18"})) inner18(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[607:592]}),({process_input[591:576]})}), .process_output(inner18_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner19"})) inner19(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[639:624]}),({process_input[623:608]})}), .process_output(inner19_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner20"})) inner20(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[671:656]}),({process_input[655:640]})}), .process_output(inner20_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner21"})) inner21(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[703:688]}),({process_input[687:672]})}), .process_output(inner21_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner22"})) inner22(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[735:720]}),({process_input[719:704]})}), .process_output(inner22_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner23"})) inner23(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[767:752]}),({process_input[751:736]})}), .process_output(inner23_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner24"})) inner24(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[799:784]}),({process_input[783:768]})}), .process_output(inner24_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner25"})) inner25(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[831:816]}),({process_input[815:800]})}), .process_output(inner25_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner26"})) inner26(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[863:848]}),({process_input[847:832]})}), .process_output(inner26_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner27"})) inner27(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[895:880]}),({process_input[879:864]})}), .process_output(inner27_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner28"})) inner28(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[927:912]}),({process_input[911:896]})}), .process_output(inner28_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner29"})) inner29(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[959:944]}),({process_input[943:928]})}), .process_output(inner29_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner30"})) inner30(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[991:976]}),({process_input[975:960]})}), .process_output(inner30_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner31"})) inner31(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1023:1008]}),({process_input[1007:992]})}), .process_output(inner31_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner32"})) inner32(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1055:1040]}),({process_input[1039:1024]})}), .process_output(inner32_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner33"})) inner33(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1087:1072]}),({process_input[1071:1056]})}), .process_output(inner33_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner34"})) inner34(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1119:1104]}),({process_input[1103:1088]})}), .process_output(inner34_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner35"})) inner35(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1151:1136]}),({process_input[1135:1120]})}), .process_output(inner35_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner36"})) inner36(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1183:1168]}),({process_input[1167:1152]})}), .process_output(inner36_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner37"})) inner37(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1215:1200]}),({process_input[1199:1184]})}), .process_output(inner37_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner38"})) inner38(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1247:1232]}),({process_input[1231:1216]})}), .process_output(inner38_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner39"})) inner39(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1279:1264]}),({process_input[1263:1248]})}), .process_output(inner39_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner40"})) inner40(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1311:1296]}),({process_input[1295:1280]})}), .process_output(inner40_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner41"})) inner41(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1343:1328]}),({process_input[1327:1312]})}), .process_output(inner41_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner42"})) inner42(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1375:1360]}),({process_input[1359:1344]})}), .process_output(inner42_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner43"})) inner43(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1407:1392]}),({process_input[1391:1376]})}), .process_output(inner43_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner44"})) inner44(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1439:1424]}),({process_input[1423:1408]})}), .process_output(inner44_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner45"})) inner45(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1471:1456]}),({process_input[1455:1440]})}), .process_output(inner45_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner46"})) inner46(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1503:1488]}),({process_input[1487:1472]})}), .process_output(inner46_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner47"})) inner47(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1535:1520]}),({process_input[1519:1504]})}), .process_output(inner47_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner48"})) inner48(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1567:1552]}),({process_input[1551:1536]})}), .process_output(inner48_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner49"})) inner49(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1599:1584]}),({process_input[1583:1568]})}), .process_output(inner49_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner50"})) inner50(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1631:1616]}),({process_input[1615:1600]})}), .process_output(inner50_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner51"})) inner51(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1663:1648]}),({process_input[1647:1632]})}), .process_output(inner51_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner52"})) inner52(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1695:1680]}),({process_input[1679:1664]})}), .process_output(inner52_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner53"})) inner53(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1727:1712]}),({process_input[1711:1696]})}), .process_output(inner53_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner54"})) inner54(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1759:1744]}),({process_input[1743:1728]})}), .process_output(inner54_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner55"})) inner55(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1791:1776]}),({process_input[1775:1760]})}), .process_output(inner55_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner56"})) inner56(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1823:1808]}),({process_input[1807:1792]})}), .process_output(inner56_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner57"})) inner57(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1855:1840]}),({process_input[1839:1824]})}), .process_output(inner57_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner58"})) inner58(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1887:1872]}),({process_input[1871:1856]})}), .process_output(inner58_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner59"})) inner59(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1919:1904]}),({process_input[1903:1888]})}), .process_output(inner59_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner60"})) inner60(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1951:1936]}),({process_input[1935:1920]})}), .process_output(inner60_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner61"})) inner61(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[1983:1968]}),({process_input[1967:1952]})}), .process_output(inner61_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner62"})) inner62(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2015:2000]}),({process_input[1999:1984]})}), .process_output(inner62_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner63"})) inner63(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2047:2032]}),({process_input[2031:2016]})}), .process_output(inner63_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner64"})) inner64(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2079:2064]}),({process_input[2063:2048]})}), .process_output(inner64_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner65"})) inner65(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2111:2096]}),({process_input[2095:2080]})}), .process_output(inner65_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner66"})) inner66(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2143:2128]}),({process_input[2127:2112]})}), .process_output(inner66_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner67"})) inner67(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2175:2160]}),({process_input[2159:2144]})}), .process_output(inner67_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner68"})) inner68(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2207:2192]}),({process_input[2191:2176]})}), .process_output(inner68_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner69"})) inner69(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2239:2224]}),({process_input[2223:2208]})}), .process_output(inner69_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner70"})) inner70(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2271:2256]}),({process_input[2255:2240]})}), .process_output(inner70_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner71"})) inner71(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2303:2288]}),({process_input[2287:2272]})}), .process_output(inner71_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner72"})) inner72(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2335:2320]}),({process_input[2319:2304]})}), .process_output(inner72_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner73"})) inner73(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2367:2352]}),({process_input[2351:2336]})}), .process_output(inner73_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner74"})) inner74(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2399:2384]}),({process_input[2383:2368]})}), .process_output(inner74_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner75"})) inner75(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2431:2416]}),({process_input[2415:2400]})}), .process_output(inner75_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner76"})) inner76(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2463:2448]}),({process_input[2447:2432]})}), .process_output(inner76_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner77"})) inner77(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2495:2480]}),({process_input[2479:2464]})}), .process_output(inner77_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner78"})) inner78(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2527:2512]}),({process_input[2511:2496]})}), .process_output(inner78_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner79"})) inner79(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2559:2544]}),({process_input[2543:2528]})}), .process_output(inner79_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner80"})) inner80(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2591:2576]}),({process_input[2575:2560]})}), .process_output(inner80_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner81"})) inner81(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2623:2608]}),({process_input[2607:2592]})}), .process_output(inner81_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner82"})) inner82(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2655:2640]}),({process_input[2639:2624]})}), .process_output(inner82_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner83"})) inner83(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2687:2672]}),({process_input[2671:2656]})}), .process_output(inner83_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner84"})) inner84(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2719:2704]}),({process_input[2703:2688]})}), .process_output(inner84_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner85"})) inner85(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2751:2736]}),({process_input[2735:2720]})}), .process_output(inner85_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner86"})) inner86(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2783:2768]}),({process_input[2767:2752]})}), .process_output(inner86_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner87"})) inner87(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2815:2800]}),({process_input[2799:2784]})}), .process_output(inner87_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner88"})) inner88(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2847:2832]}),({process_input[2831:2816]})}), .process_output(inner88_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner89"})) inner89(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2879:2864]}),({process_input[2863:2848]})}), .process_output(inner89_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner90"})) inner90(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2911:2896]}),({process_input[2895:2880]})}), .process_output(inner90_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner91"})) inner91(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2943:2928]}),({process_input[2927:2912]})}), .process_output(inner91_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner92"})) inner92(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[2975:2960]}),({process_input[2959:2944]})}), .process_output(inner92_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner93"})) inner93(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3007:2992]}),({process_input[2991:2976]})}), .process_output(inner93_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner94"})) inner94(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3039:3024]}),({process_input[3023:3008]})}), .process_output(inner94_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner95"})) inner95(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3071:3056]}),({process_input[3055:3040]})}), .process_output(inner95_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner96"})) inner96(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3103:3088]}),({process_input[3087:3072]})}), .process_output(inner96_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner97"})) inner97(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3135:3120]}),({process_input[3119:3104]})}), .process_output(inner97_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner98"})) inner98(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3167:3152]}),({process_input[3151:3136]})}), .process_output(inner98_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner99"})) inner99(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3199:3184]}),({process_input[3183:3168]})}), .process_output(inner99_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner100"})) inner100(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3231:3216]}),({process_input[3215:3200]})}), .process_output(inner100_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner101"})) inner101(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3263:3248]}),({process_input[3247:3232]})}), .process_output(inner101_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner102"})) inner102(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3295:3280]}),({process_input[3279:3264]})}), .process_output(inner102_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner103"})) inner103(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3327:3312]}),({process_input[3311:3296]})}), .process_output(inner103_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner104"})) inner104(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3359:3344]}),({process_input[3343:3328]})}), .process_output(inner104_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner105"})) inner105(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3391:3376]}),({process_input[3375:3360]})}), .process_output(inner105_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner106"})) inner106(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3423:3408]}),({process_input[3407:3392]})}), .process_output(inner106_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner107"})) inner107(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3455:3440]}),({process_input[3439:3424]})}), .process_output(inner107_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner108"})) inner108(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3487:3472]}),({process_input[3471:3456]})}), .process_output(inner108_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner109"})) inner109(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3519:3504]}),({process_input[3503:3488]})}), .process_output(inner109_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner110"})) inner110(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3551:3536]}),({process_input[3535:3520]})}), .process_output(inner110_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner111"})) inner111(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3583:3568]}),({process_input[3567:3552]})}), .process_output(inner111_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner112"})) inner112(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3615:3600]}),({process_input[3599:3584]})}), .process_output(inner112_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner113"})) inner113(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3647:3632]}),({process_input[3631:3616]})}), .process_output(inner113_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner114"})) inner114(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3679:3664]}),({process_input[3663:3648]})}), .process_output(inner114_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner115"})) inner115(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3711:3696]}),({process_input[3695:3680]})}), .process_output(inner115_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner116"})) inner116(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3743:3728]}),({process_input[3727:3712]})}), .process_output(inner116_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner117"})) inner117(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3775:3760]}),({process_input[3759:3744]})}), .process_output(inner117_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner118"})) inner118(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3807:3792]}),({process_input[3791:3776]})}), .process_output(inner118_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner119"})) inner119(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3839:3824]}),({process_input[3823:3808]})}), .process_output(inner119_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner120"})) inner120(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3871:3856]}),({process_input[3855:3840]})}), .process_output(inner120_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner121"})) inner121(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3903:3888]}),({process_input[3887:3872]})}), .process_output(inner121_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner122"})) inner122(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3935:3920]}),({process_input[3919:3904]})}), .process_output(inner122_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner123"})) inner123(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3967:3952]}),({process_input[3951:3936]})}), .process_output(inner123_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner124"})) inner124(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[3999:3984]}),({process_input[3983:3968]})}), .process_output(inner124_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner125"})) inner125(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[4031:4016]}),({process_input[4015:4000]})}), .process_output(inner125_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner126"})) inner126(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[4063:4048]}),({process_input[4047:4032]})}), .process_output(inner126_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner127"})) inner127(.CLK(CLK), .process_CE(process_CE), .sum_inp({({process_input[4095:4080]}),({process_input[4079:4064]})}), .process_output(inner127_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner128"})) inner128(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner1_process_output,inner0_process_output}), .process_output(inner128_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner129"})) inner129(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner3_process_output,inner2_process_output}), .process_output(inner129_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner130"})) inner130(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner5_process_output,inner4_process_output}), .process_output(inner130_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner131"})) inner131(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner7_process_output,inner6_process_output}), .process_output(inner131_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner132"})) inner132(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner9_process_output,inner8_process_output}), .process_output(inner132_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner133"})) inner133(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner11_process_output,inner10_process_output}), .process_output(inner133_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner134"})) inner134(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner13_process_output,inner12_process_output}), .process_output(inner134_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner135"})) inner135(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner15_process_output,inner14_process_output}), .process_output(inner135_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner136"})) inner136(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner17_process_output,inner16_process_output}), .process_output(inner136_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner137"})) inner137(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner19_process_output,inner18_process_output}), .process_output(inner137_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner138"})) inner138(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner21_process_output,inner20_process_output}), .process_output(inner138_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner139"})) inner139(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner23_process_output,inner22_process_output}), .process_output(inner139_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner140"})) inner140(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner25_process_output,inner24_process_output}), .process_output(inner140_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner141"})) inner141(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner27_process_output,inner26_process_output}), .process_output(inner141_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner142"})) inner142(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner29_process_output,inner28_process_output}), .process_output(inner142_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner143"})) inner143(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner31_process_output,inner30_process_output}), .process_output(inner143_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner144"})) inner144(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner33_process_output,inner32_process_output}), .process_output(inner144_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner145"})) inner145(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner35_process_output,inner34_process_output}), .process_output(inner145_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner146"})) inner146(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner37_process_output,inner36_process_output}), .process_output(inner146_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner147"})) inner147(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner39_process_output,inner38_process_output}), .process_output(inner147_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner148"})) inner148(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner41_process_output,inner40_process_output}), .process_output(inner148_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner149"})) inner149(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner43_process_output,inner42_process_output}), .process_output(inner149_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner150"})) inner150(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner45_process_output,inner44_process_output}), .process_output(inner150_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner151"})) inner151(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner47_process_output,inner46_process_output}), .process_output(inner151_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner152"})) inner152(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner49_process_output,inner48_process_output}), .process_output(inner152_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner153"})) inner153(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner51_process_output,inner50_process_output}), .process_output(inner153_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner154"})) inner154(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner53_process_output,inner52_process_output}), .process_output(inner154_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner155"})) inner155(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner55_process_output,inner54_process_output}), .process_output(inner155_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner156"})) inner156(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner57_process_output,inner56_process_output}), .process_output(inner156_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner157"})) inner157(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner59_process_output,inner58_process_output}), .process_output(inner157_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner158"})) inner158(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner61_process_output,inner60_process_output}), .process_output(inner158_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner159"})) inner159(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner63_process_output,inner62_process_output}), .process_output(inner159_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner160"})) inner160(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner65_process_output,inner64_process_output}), .process_output(inner160_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner161"})) inner161(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner67_process_output,inner66_process_output}), .process_output(inner161_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner162"})) inner162(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner69_process_output,inner68_process_output}), .process_output(inner162_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner163"})) inner163(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner71_process_output,inner70_process_output}), .process_output(inner163_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner164"})) inner164(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner73_process_output,inner72_process_output}), .process_output(inner164_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner165"})) inner165(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner75_process_output,inner74_process_output}), .process_output(inner165_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner166"})) inner166(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner77_process_output,inner76_process_output}), .process_output(inner166_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner167"})) inner167(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner79_process_output,inner78_process_output}), .process_output(inner167_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner168"})) inner168(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner81_process_output,inner80_process_output}), .process_output(inner168_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner169"})) inner169(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner83_process_output,inner82_process_output}), .process_output(inner169_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner170"})) inner170(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner85_process_output,inner84_process_output}), .process_output(inner170_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner171"})) inner171(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner87_process_output,inner86_process_output}), .process_output(inner171_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner172"})) inner172(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner89_process_output,inner88_process_output}), .process_output(inner172_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner173"})) inner173(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner91_process_output,inner90_process_output}), .process_output(inner173_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner174"})) inner174(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner93_process_output,inner92_process_output}), .process_output(inner174_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner175"})) inner175(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner95_process_output,inner94_process_output}), .process_output(inner175_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner176"})) inner176(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner97_process_output,inner96_process_output}), .process_output(inner176_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner177"})) inner177(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner99_process_output,inner98_process_output}), .process_output(inner177_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner178"})) inner178(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner101_process_output,inner100_process_output}), .process_output(inner178_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner179"})) inner179(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner103_process_output,inner102_process_output}), .process_output(inner179_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner180"})) inner180(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner105_process_output,inner104_process_output}), .process_output(inner180_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner181"})) inner181(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner107_process_output,inner106_process_output}), .process_output(inner181_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner182"})) inner182(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner109_process_output,inner108_process_output}), .process_output(inner182_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner183"})) inner183(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner111_process_output,inner110_process_output}), .process_output(inner183_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner184"})) inner184(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner113_process_output,inner112_process_output}), .process_output(inner184_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner185"})) inner185(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner115_process_output,inner114_process_output}), .process_output(inner185_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner186"})) inner186(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner117_process_output,inner116_process_output}), .process_output(inner186_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner187"})) inner187(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner119_process_output,inner118_process_output}), .process_output(inner187_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner188"})) inner188(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner121_process_output,inner120_process_output}), .process_output(inner188_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner189"})) inner189(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner123_process_output,inner122_process_output}), .process_output(inner189_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner190"})) inner190(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner125_process_output,inner124_process_output}), .process_output(inner190_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner191"})) inner191(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner127_process_output,inner126_process_output}), .process_output(inner191_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner192"})) inner192(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner129_process_output,inner128_process_output}), .process_output(inner192_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner193"})) inner193(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner131_process_output,inner130_process_output}), .process_output(inner193_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner194"})) inner194(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner133_process_output,inner132_process_output}), .process_output(inner194_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner195"})) inner195(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner135_process_output,inner134_process_output}), .process_output(inner195_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner196"})) inner196(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner137_process_output,inner136_process_output}), .process_output(inner196_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner197"})) inner197(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner139_process_output,inner138_process_output}), .process_output(inner197_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner198"})) inner198(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner141_process_output,inner140_process_output}), .process_output(inner198_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner199"})) inner199(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner143_process_output,inner142_process_output}), .process_output(inner199_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner200"})) inner200(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner145_process_output,inner144_process_output}), .process_output(inner200_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner201"})) inner201(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner147_process_output,inner146_process_output}), .process_output(inner201_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner202"})) inner202(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner149_process_output,inner148_process_output}), .process_output(inner202_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner203"})) inner203(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner151_process_output,inner150_process_output}), .process_output(inner203_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner204"})) inner204(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner153_process_output,inner152_process_output}), .process_output(inner204_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner205"})) inner205(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner155_process_output,inner154_process_output}), .process_output(inner205_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner206"})) inner206(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner157_process_output,inner156_process_output}), .process_output(inner206_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner207"})) inner207(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner159_process_output,inner158_process_output}), .process_output(inner207_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner208"})) inner208(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner161_process_output,inner160_process_output}), .process_output(inner208_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner209"})) inner209(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner163_process_output,inner162_process_output}), .process_output(inner209_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner210"})) inner210(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner165_process_output,inner164_process_output}), .process_output(inner210_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner211"})) inner211(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner167_process_output,inner166_process_output}), .process_output(inner211_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner212"})) inner212(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner169_process_output,inner168_process_output}), .process_output(inner212_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner213"})) inner213(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner171_process_output,inner170_process_output}), .process_output(inner213_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner214"})) inner214(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner173_process_output,inner172_process_output}), .process_output(inner214_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner215"})) inner215(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner175_process_output,inner174_process_output}), .process_output(inner215_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner216"})) inner216(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner177_process_output,inner176_process_output}), .process_output(inner216_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner217"})) inner217(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner179_process_output,inner178_process_output}), .process_output(inner217_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner218"})) inner218(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner181_process_output,inner180_process_output}), .process_output(inner218_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner219"})) inner219(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner183_process_output,inner182_process_output}), .process_output(inner219_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner220"})) inner220(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner185_process_output,inner184_process_output}), .process_output(inner220_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner221"})) inner221(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner187_process_output,inner186_process_output}), .process_output(inner221_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner222"})) inner222(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner189_process_output,inner188_process_output}), .process_output(inner222_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner223"})) inner223(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner191_process_output,inner190_process_output}), .process_output(inner223_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner224"})) inner224(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner193_process_output,inner192_process_output}), .process_output(inner224_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner225"})) inner225(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner195_process_output,inner194_process_output}), .process_output(inner225_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner226"})) inner226(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner197_process_output,inner196_process_output}), .process_output(inner226_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner227"})) inner227(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner199_process_output,inner198_process_output}), .process_output(inner227_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner228"})) inner228(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner201_process_output,inner200_process_output}), .process_output(inner228_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner229"})) inner229(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner203_process_output,inner202_process_output}), .process_output(inner229_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner230"})) inner230(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner205_process_output,inner204_process_output}), .process_output(inner230_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner231"})) inner231(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner207_process_output,inner206_process_output}), .process_output(inner231_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner232"})) inner232(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner209_process_output,inner208_process_output}), .process_output(inner232_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner233"})) inner233(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner211_process_output,inner210_process_output}), .process_output(inner233_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner234"})) inner234(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner213_process_output,inner212_process_output}), .process_output(inner234_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner235"})) inner235(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner215_process_output,inner214_process_output}), .process_output(inner235_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner236"})) inner236(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner217_process_output,inner216_process_output}), .process_output(inner236_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner237"})) inner237(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner219_process_output,inner218_process_output}), .process_output(inner237_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner238"})) inner238(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner221_process_output,inner220_process_output}), .process_output(inner238_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner239"})) inner239(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner223_process_output,inner222_process_output}), .process_output(inner239_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner240"})) inner240(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner225_process_output,inner224_process_output}), .process_output(inner240_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner241"})) inner241(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner227_process_output,inner226_process_output}), .process_output(inner241_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner242"})) inner242(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner229_process_output,inner228_process_output}), .process_output(inner242_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner243"})) inner243(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner231_process_output,inner230_process_output}), .process_output(inner243_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner244"})) inner244(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner233_process_output,inner232_process_output}), .process_output(inner244_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner245"})) inner245(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner235_process_output,inner234_process_output}), .process_output(inner245_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner246"})) inner246(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner237_process_output,inner236_process_output}), .process_output(inner246_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner247"})) inner247(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner239_process_output,inner238_process_output}), .process_output(inner247_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner248"})) inner248(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner241_process_output,inner240_process_output}), .process_output(inner248_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner249"})) inner249(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner243_process_output,inner242_process_output}), .process_output(inner249_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner250"})) inner250(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner245_process_output,inner244_process_output}), .process_output(inner250_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner251"})) inner251(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner247_process_output,inner246_process_output}), .process_output(inner251_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner252"})) inner252(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner249_process_output,inner248_process_output}), .process_output(inner252_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner253"})) inner253(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner251_process_output,inner250_process_output}), .process_output(inner253_process_output));
  ABS_SUM #(.INSTANCE_NAME({INSTANCE_NAME,"_inner254"})) inner254(.CLK(CLK), .process_CE(process_CE), .sum_inp({inner253_process_output,inner252_process_output}), .process_output(inner254_process_output));
endmodule

module SAD(input CLK, input CE, input [4095:0] process_input, output [15:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [4095:0] partial_process_output;
  wire [15:0] sum_process_output;
  assign process_output = sum_process_output;
  // function: process pure=true delay=11
  // function: reset pure=true delay=0
  map_absoluteDiff_W16_H16 #(.INSTANCE_NAME({INSTANCE_NAME,"_partial"})) partial(.CLK(CLK), .process_CE(CE), .process_input(process_input), .process_output(partial_process_output));
  reduce_ABS_SUM_W16_H16 #(.INSTANCE_NAME({INSTANCE_NAME,"_sum"})) sum(.CLK(CLK), .process_CE(CE), .process_input(partial_process_output), .process_output(sum_process_output));
endmodule

module map_SAD_W2_H1(input CLK, input process_CE, input [8191:0] process_input, output [31:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] inner0_0_process_output;
  wire [15:0] inner1_0_process_output;
  assign process_output = {inner1_0_process_output,inner0_0_process_output};
  // function: process pure=true delay=11
  SAD #(.INSTANCE_NAME({INSTANCE_NAME,"_inner0_0"})) inner0_0(.CLK(CLK), .CE(process_CE), .process_input(({process_input[4095:0]})), .process_output(inner0_0_process_output));
  SAD #(.INSTANCE_NAME({INSTANCE_NAME,"_inner1_0"})) inner1_0(.CLK(CLK), .CE(process_CE), .process_input(({process_input[8191:4096]})), .process_output(inner1_0_process_output));
endmodule

module LowerSum(input CLK, input process_CE, input [15:0] LOWER_SUM_INP, output [15:0] process_output);
parameter INSTANCE_NAME="INST";
  assign process_output = LOWER_SUM_INP;
  // function: process pure=true delay=0
endmodule

module map_LowerSum_W2_H1(input CLK, input process_CE, input [31:0] process_input, output [31:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] inner0_0_process_output;
  wire [15:0] inner1_0_process_output;
  assign process_output = {inner1_0_process_output,inner0_0_process_output};
  // function: process pure=true delay=0
  LowerSum #(.INSTANCE_NAME({INSTANCE_NAME,"_inner0_0"})) inner0_0(.CLK(CLK), .process_CE(process_CE), .LOWER_SUM_INP(({process_input[15:0]})), .process_output(inner0_0_process_output));
  LowerSum #(.INSTANCE_NAME({INSTANCE_NAME,"_inner1_0"})) inner1_0(.CLK(CLK), .process_CE(process_CE), .LOWER_SUM_INP(({process_input[31:16]})), .process_output(inner1_0_process_output));
endmodule

module packTupleArrays_table__0x470eb890(input CLK, input process_CE, input [47:0] process_input, output [47:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [15:0] unnamedcast34551USEDMULTIPLEcast;assign unnamedcast34551USEDMULTIPLEcast = (process_input[15:0]); 
  wire [31:0] unnamedcast34555USEDMULTIPLEcast;assign unnamedcast34555USEDMULTIPLEcast = (process_input[47:16]); 
  assign process_output = {{({unnamedcast34555USEDMULTIPLEcast[31:16]}),({unnamedcast34551USEDMULTIPLEcast[15:8]})},{({unnamedcast34555USEDMULTIPLEcast[15:0]}),({unnamedcast34551USEDMULTIPLEcast[7:0]})}};
  // function: process pure=true delay=0
endmodule

module argmin_asyncnil(input CLK, input process_CE, input [47:0] inp, output [23:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [23:0] unnamedcast34571USEDMULTIPLEcast;assign unnamedcast34571USEDMULTIPLEcast = (inp[23:0]); 
  wire [23:0] unnamedcast34575USEDMULTIPLEcast;assign unnamedcast34575USEDMULTIPLEcast = (inp[47:24]); 
  reg unnamedbinop34578_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedbinop34578_delay1_validunnamednull0_CEprocess_CE <= {(((unnamedcast34571USEDMULTIPLEcast[23:8]))<=((unnamedcast34575USEDMULTIPLEcast[23:8])))}; end end
  reg [23:0] unnamedcast34571_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast34571_delay1_validunnamednull0_CEprocess_CE <= unnamedcast34571USEDMULTIPLEcast; end end
  reg [23:0] unnamedcast34575_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedcast34575_delay1_validunnamednull0_CEprocess_CE <= unnamedcast34575USEDMULTIPLEcast; end end
  reg [23:0] unnamedselect34579_delay1_validunnamednull0_CEprocess_CE;  always @ (posedge CLK) begin if (process_CE) begin unnamedselect34579_delay1_validunnamednull0_CEprocess_CE <= ((unnamedbinop34578_delay1_validunnamednull0_CEprocess_CE)?(unnamedcast34571_delay1_validunnamednull0_CEprocess_CE):(unnamedcast34575_delay1_validunnamednull0_CEprocess_CE)); end end
  assign process_output = unnamedselect34579_delay1_validunnamednull0_CEprocess_CE;
  // function: process pure=true delay=2
endmodule

module reduce_argmin_asyncnil_W2_H1(input CLK, input process_CE, input [47:0] process_input, output [23:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [23:0] inner0_process_output;
  assign process_output = inner0_process_output;
  // function: process pure=true delay=2
  argmin_asyncnil #(.INSTANCE_NAME({INSTANCE_NAME,"_inner0"})) inner0(.CLK(CLK), .process_CE(process_CE), .inp({({process_input[47:24]}),({process_input[23:0]})}), .process_output(inner0_process_output));
endmodule

module argmin_asynctrue(input CLK, input process_CE, input [47:0] inp, output [23:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [23:0] unnamedcast34601USEDMULTIPLEcast;assign unnamedcast34601USEDMULTIPLEcast = (inp[23:0]); 
  wire [23:0] unnamedcast34605USEDMULTIPLEcast;assign unnamedcast34605USEDMULTIPLEcast = (inp[47:24]); 
  assign process_output = (({(((unnamedcast34601USEDMULTIPLEcast[23:8]))<=((unnamedcast34605USEDMULTIPLEcast[23:8])))})?(unnamedcast34601USEDMULTIPLEcast):(unnamedcast34605USEDMULTIPLEcast));
  // function: process pure=true delay=0
endmodule

module RegBy_argmin_asynctrue_CEtrue_initnil(input CLK, input set_valid, input CE, input [23:0] set_inp, input setby_valid, input [23:0] setby_inp, output [23:0] SETBY_OUTPUT, output [23:0] GET_OUTPUT);
parameter INSTANCE_NAME="INST";
  reg [23:0] R;
  wire [23:0] regby_inner_process_output;
  always @(posedge CLK) begin if(set_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(setby_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,set_valid})+({4'b0,setby_valid})) > 5'd1) begin $display("error, function 'set' on instance 'R' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [24:0] unnamedcallArbitrate34644USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate34644USEDMULTIPLEcallArbitrate = {(set_valid||setby_valid),((set_valid)?(set_inp):(regby_inner_process_output))}; 
    always @ (posedge CLK) begin if ((unnamedcallArbitrate34644USEDMULTIPLEcallArbitrate[24]) && CE) begin R <= (unnamedcallArbitrate34644USEDMULTIPLEcallArbitrate[23:0]); end end
  assign SETBY_OUTPUT = regby_inner_process_output;
  assign GET_OUTPUT = R;
  // function: set pure=false ONLY WIRE
  // function: setby pure=false ONLY WIRE
  // function: get pure=true ONLY WIRE
  argmin_asynctrue #(.INSTANCE_NAME({INSTANCE_NAME,"_regby_inner"})) regby_inner(.CLK(CLK), .process_CE(CE), .inp({setby_inp,R}), .process_output(regby_inner_process_output));
endmodule

module ReduceSeq_argmin_asynctrue_T8(input CLK, input process_valid, input CE, input [23:0] process_input, output [24:0] process_output, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  wire [15:0] phase_GET_OUTPUT;
  wire unnamedbinop34658USEDMULTIPLEbinop;assign unnamedbinop34658USEDMULTIPLEbinop = {(phase_GET_OUTPUT==(16'd0))}; 
  wire [23:0] result_SETBY_OUTPUT;
  reg [23:0] unnamedcall34660_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcall34660_delay1_validunnamednull0_CECE <= result_SETBY_OUTPUT; end end
  reg unnamedbinop34664_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedbinop34664_delay1_validunnamednull0_CECE <= {(phase_GET_OUTPUT==(16'd7))}; end end
  wire [15:0] phase_SETBY_OUTPUT;
  assign process_output = {unnamedbinop34664_delay1_validunnamednull0_CECE,unnamedcall34660_delay1_validunnamednull0_CECE};
  // function: process pure=false delay=1
  // function: reset pure=false delay=0
  RegBy_sumwrap_uint16_to7_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_phase"})) phase(.CLK(CLK), .set_valid(reset), .CE(CE), .set_inp((16'd0)), .setby_valid(process_valid), .setby_inp((16'd1)), .SETBY_OUTPUT(phase_SETBY_OUTPUT), .GET_OUTPUT(phase_GET_OUTPUT));
  RegBy_argmin_asynctrue_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_result"})) result(.CLK(CLK), .set_valid({(unnamedbinop34658USEDMULTIPLEbinop&&process_valid)}), .CE(CE), .set_inp(process_input), .setby_valid({({(~unnamedbinop34658USEDMULTIPLEbinop)}&&process_valid)}), .setby_inp(process_input), .SETBY_OUTPUT(result_SETBY_OUTPUT), .GET_OUTPUT(result_GET_OUTPUT));
endmodule

module argmin(input CLK, input process_valid, input CE, input [8191:0] process_input, output [24:0] process_output, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  wire [15:0] convKernel_process_output;
  reg [15:0] unnamedcall34706_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcall34706_delay1_validunnamednull0_CECE <= convKernel_process_output; end end
  reg [15:0] unnamedcall34706_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcall34706_delay2_validunnamednull0_CECE <= unnamedcall34706_delay1_validunnamednull0_CECE; end end
  reg [15:0] unnamedcall34706_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcall34706_delay3_validunnamednull0_CECE <= unnamedcall34706_delay2_validunnamednull0_CECE; end end
  reg [15:0] unnamedcall34706_delay4_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcall34706_delay4_validunnamednull0_CECE <= unnamedcall34706_delay3_validunnamednull0_CECE; end end
  reg [15:0] unnamedcall34706_delay5_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcall34706_delay5_validunnamednull0_CECE <= unnamedcall34706_delay4_validunnamednull0_CECE; end end
  reg [15:0] unnamedcall34706_delay6_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcall34706_delay6_validunnamednull0_CECE <= unnamedcall34706_delay5_validunnamednull0_CECE; end end
  reg [15:0] unnamedcall34706_delay7_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcall34706_delay7_validunnamednull0_CECE <= unnamedcall34706_delay6_validunnamednull0_CECE; end end
  reg [15:0] unnamedcall34706_delay8_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcall34706_delay8_validunnamednull0_CECE <= unnamedcall34706_delay7_validunnamednull0_CECE; end end
  reg [15:0] unnamedcall34706_delay9_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcall34706_delay9_validunnamednull0_CECE <= unnamedcall34706_delay8_validunnamednull0_CECE; end end
  reg [15:0] unnamedcall34706_delay10_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcall34706_delay10_validunnamednull0_CECE <= unnamedcall34706_delay9_validunnamednull0_CECE; end end
  reg [15:0] unnamedcall34706_delay11_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcall34706_delay11_validunnamednull0_CECE <= unnamedcall34706_delay10_validunnamednull0_CECE; end end
  wire [31:0] sadvalues_process_output;
  wire [31:0] LOWER_SUM_process_output;
  wire [47:0] SOS_process_output;
  wire [23:0] argmin_process_output;
  reg process_valid_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay1_validunnamednull0_CECE <= process_valid; end end
  reg process_valid_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay2_validunnamednull0_CECE <= process_valid_delay1_validunnamednull0_CECE; end end
  reg process_valid_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay3_validunnamednull0_CECE <= process_valid_delay2_validunnamednull0_CECE; end end
  reg process_valid_delay4_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay4_validunnamednull0_CECE <= process_valid_delay3_validunnamednull0_CECE; end end
  reg process_valid_delay5_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay5_validunnamednull0_CECE <= process_valid_delay4_validunnamednull0_CECE; end end
  reg process_valid_delay6_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay6_validunnamednull0_CECE <= process_valid_delay5_validunnamednull0_CECE; end end
  reg process_valid_delay7_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay7_validunnamednull0_CECE <= process_valid_delay6_validunnamednull0_CECE; end end
  reg process_valid_delay8_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay8_validunnamednull0_CECE <= process_valid_delay7_validunnamednull0_CECE; end end
  reg process_valid_delay9_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay9_validunnamednull0_CECE <= process_valid_delay8_validunnamednull0_CECE; end end
  reg process_valid_delay10_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay10_validunnamednull0_CECE <= process_valid_delay9_validunnamednull0_CECE; end end
  reg process_valid_delay11_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay11_validunnamednull0_CECE <= process_valid_delay10_validunnamednull0_CECE; end end
  reg process_valid_delay12_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay12_validunnamednull0_CECE <= process_valid_delay11_validunnamednull0_CECE; end end
  reg process_valid_delay13_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_valid_delay13_validunnamednull0_CECE <= process_valid_delay12_validunnamednull0_CECE; end end
  wire [24:0] argminseq_process_output;
  assign process_output = argminseq_process_output;
  // function: process pure=false delay=14
  // function: reset pure=false delay=0
  constSeq_table__0x44c9de70_T8 #(.INSTANCE_NAME({INSTANCE_NAME,"_convKernel"})) convKernel(.CLK(CLK), .process_valid(process_valid), .process_CE(CE), .process_output(convKernel_process_output));
  map_SAD_W2_H1 #(.INSTANCE_NAME({INSTANCE_NAME,"_sadvalues"})) sadvalues(.CLK(CLK), .process_CE(CE), .process_input(process_input), .process_output(sadvalues_process_output));
  map_LowerSum_W2_H1 #(.INSTANCE_NAME({INSTANCE_NAME,"_LOWER_SUM"})) LOWER_SUM(.CLK(CLK), .process_CE(CE), .process_input(sadvalues_process_output), .process_output(LOWER_SUM_process_output));
  packTupleArrays_table__0x470eb890 #(.INSTANCE_NAME({INSTANCE_NAME,"_SOS"})) SOS(.CLK(CLK), .process_CE(CE), .process_input({LOWER_SUM_process_output,unnamedcall34706_delay11_validunnamednull0_CECE}), .process_output(SOS_process_output));
  reduce_argmin_asyncnil_W2_H1 #(.INSTANCE_NAME({INSTANCE_NAME,"_argmin"})) argmin(.CLK(CLK), .process_CE(CE), .process_input(SOS_process_output), .process_output(argmin_process_output));
  ReduceSeq_argmin_asynctrue_T8 #(.INSTANCE_NAME({INSTANCE_NAME,"_argminseq"})) argminseq(.CLK(CLK), .process_valid(process_valid_delay13_validunnamednull0_CECE), .CE(CE), .process_input(argmin_process_output), .process_output(argminseq_process_output), .reset(reset));
endmodule

module LiftDecimate_argmin(input CLK, output ready, input reset, input CE, input process_valid, input [8192:0] process_input, output [24:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  assign ready = (1'd1);
  wire unnamedcast34880USEDMULTIPLEcast;assign unnamedcast34880USEDMULTIPLEcast = (process_input[8192]); 
  wire [24:0] LiftDecimate_process_output;
  reg [23:0] unnamedcast34883_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast34883_delay1_validunnamednull0_CECE <= (LiftDecimate_process_output[23:0]); end end
  reg unnamedcast34880_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast34880_delay1_validunnamednull0_CECE <= unnamedcast34880USEDMULTIPLEcast; end end
  reg unnamedcast34880_delay2_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast34880_delay2_validunnamednull0_CECE <= unnamedcast34880_delay1_validunnamednull0_CECE; end end
  reg unnamedcast34880_delay3_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast34880_delay3_validunnamednull0_CECE <= unnamedcast34880_delay2_validunnamednull0_CECE; end end
  reg unnamedcast34880_delay4_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast34880_delay4_validunnamednull0_CECE <= unnamedcast34880_delay3_validunnamednull0_CECE; end end
  reg unnamedcast34880_delay5_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast34880_delay5_validunnamednull0_CECE <= unnamedcast34880_delay4_validunnamednull0_CECE; end end
  reg unnamedcast34880_delay6_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast34880_delay6_validunnamednull0_CECE <= unnamedcast34880_delay5_validunnamednull0_CECE; end end
  reg unnamedcast34880_delay7_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast34880_delay7_validunnamednull0_CECE <= unnamedcast34880_delay6_validunnamednull0_CECE; end end
  reg unnamedcast34880_delay8_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast34880_delay8_validunnamednull0_CECE <= unnamedcast34880_delay7_validunnamednull0_CECE; end end
  reg unnamedcast34880_delay9_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast34880_delay9_validunnamednull0_CECE <= unnamedcast34880_delay8_validunnamednull0_CECE; end end
  reg unnamedcast34880_delay10_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast34880_delay10_validunnamednull0_CECE <= unnamedcast34880_delay9_validunnamednull0_CECE; end end
  reg unnamedcast34880_delay11_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast34880_delay11_validunnamednull0_CECE <= unnamedcast34880_delay10_validunnamednull0_CECE; end end
  reg unnamedcast34880_delay12_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast34880_delay12_validunnamednull0_CECE <= unnamedcast34880_delay11_validunnamednull0_CECE; end end
  reg unnamedcast34880_delay13_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast34880_delay13_validunnamednull0_CECE <= unnamedcast34880_delay12_validunnamednull0_CECE; end end
  reg unnamedcast34880_delay14_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast34880_delay14_validunnamednull0_CECE <= unnamedcast34880_delay13_validunnamednull0_CECE; end end
  reg unnamedbinop34888_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedbinop34888_delay1_validunnamednull0_CECE <= {((LiftDecimate_process_output[24])&&unnamedcast34880_delay14_validunnamednull0_CECE)}; end end
  assign process_output = {unnamedbinop34888_delay1_validunnamednull0_CECE,unnamedcast34883_delay1_validunnamednull0_CECE};
  // function: ready pure=true delay=0
  // function: reset pure=false delay=0
  // function: process pure=false delay=15
  argmin #(.INSTANCE_NAME({INSTANCE_NAME,"_LiftDecimate"})) LiftDecimate(.CLK(CLK), .process_valid({(unnamedcast34880USEDMULTIPLEcast&&process_valid)}), .CE(CE), .process_input((process_input[8191:0])), .process_output(LiftDecimate_process_output), .reset(reset));
endmodule

module LiftHandshake_LiftDecimate_argmin(input CLK, input ready_downstream, output ready, input reset, input [8192:0] process_input, output [24:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire inner_LiftDecimate_argmin_ready;
  assign ready = {(inner_LiftDecimate_argmin_ready&&ready_downstream)};
  wire unnamedbinop34938USEDMULTIPLEbinop;assign unnamedbinop34938USEDMULTIPLEbinop = {(reset||ready_downstream)}; 
  wire unnamedunary34939USEDMULTIPLEunary;assign unnamedunary34939USEDMULTIPLEunary = {(~reset)}; 
  wire [24:0] inner_LiftDecimate_argmin_process_output;
  wire validBitDelay_LiftDecimate_argmin_pushPop_out;
  wire [24:0] unnamedtuple34949USEDMULTIPLEtuple;assign unnamedtuple34949USEDMULTIPLEtuple = {{((inner_LiftDecimate_argmin_process_output[24])&&validBitDelay_LiftDecimate_argmin_pushPop_out)},(inner_LiftDecimate_argmin_process_output[23:0])}; 
  always @(posedge CLK) begin if({(~{((unnamedtuple34949USEDMULTIPLEtuple[24])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: output valid bit should not be X!",INSTANCE_NAME); end end
  always @(posedge CLK) begin if({(~{((process_input[8192])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = unnamedtuple34949USEDMULTIPLEtuple;
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  LiftDecimate_argmin #(.INSTANCE_NAME({INSTANCE_NAME,"_inner_LiftDecimate_argmin"})) inner_LiftDecimate_argmin(.CLK(CLK), .ready(inner_LiftDecimate_argmin_ready), .reset(reset), .CE(unnamedbinop34938USEDMULTIPLEbinop), .process_valid(unnamedunary34939USEDMULTIPLEunary), .process_input(process_input), .process_output(inner_LiftDecimate_argmin_process_output));
  ShiftRegister_15_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_validBitDelay_LiftDecimate_argmin"})) validBitDelay_LiftDecimate_argmin(.CLK(CLK), .pushPop_valid(unnamedunary34939USEDMULTIPLEunary), .CE(unnamedbinop34938USEDMULTIPLEbinop), .sr_input((1'd1)), .pushPop_out(validBitDelay_LiftDecimate_argmin_pushPop_out), .reset(reset));
endmodule

module hsfn(input CLK, input ready_downstream, output ready, input reset, input [64:0] process_input, output [64:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire [3:0] unnamedtuple36533USEDMULTIPLEtuple;assign unnamedtuple36533USEDMULTIPLEtuple = {(1'd1),(1'd1),(1'd1),ready_downstream}; 
  wire f1_store_ready;
  wire left_ready;
  wire f2_store_ready;
  wire right_ready;
  wire inp_broadcast_ready;
  wire oi0_ready;
  wire pad_ready;
  wire reducerate_ready;
  wire f3_store_ready;
  wire AM_ready;
  wire mer_ready;
  wire [1:0] merge_ready;
  wire rb2_ready;
  wire right2_ready;
  wire rup_ready;
  wire rAO_ready;
  wire rightLB_ready;
  wire AOr_ready;
  wire f2_load_ready;
  wire llb_ready;
  wire LB_ready;
  wire AO_ready;
  wire f1_load_ready;
  wire incrate_ready;
  wire CRP_ready;
  wire display_ready;
  wire f3_load_ready;
  assign ready = reducerate_ready;
  wire [0:0] unnamedtuple36395USEDMULTIPLEtuple;assign unnamedtuple36395USEDMULTIPLEtuple = {(1'd1)}; 
  wire [24:0] f3_load_output;
  wire [32:0] display_process_output;
  wire [32:0] CRP_process_output;
  wire [64:0] incrate_process_output;
  wire [16:0] reducerate_process_output;
  wire [16:0] pad_process_output;
  wire [16:0] oi0_process_output;
  wire [33:0] inp_broadcast_process_output;
  wire [8:0] left_process_output;
  wire [0:0] f1_store_output;
  wire [8:0] right_process_output;
  wire [0:0] f2_store_output;
  wire [8:0] f1_load_output;
  wire [8:0] AO_process_output;
  wire [2176:0] LB_process_output;
  wire [4096:0] llb_process_output;
  wire [8:0] f2_load_output;
  wire [8:0] AOr_process_output;
  wire [2048:0] rightLB_process_output;
  wire [2048:0] rAO_process_output;
  wire [2048:0] rup_process_output;
  wire [2048:0] right2_process_output;
  wire [4096:0] rb2_process_output;
  wire [8192:0] merge_process_output;
  wire [8192:0] mer_process_output;
  wire [24:0] AM_process_output;
  wire [0:0] f3_store_output;
  assign process_output = incrate_process_output;
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  LiftHandshake_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128 #(.INSTANCE_NAME({INSTANCE_NAME,"_f1"})) f1(.CLK(CLK), .load_input(unnamedtuple36395USEDMULTIPLEtuple), .load_output(f1_load_output), .store_reset(reset), .store_ready_downstream((unnamedtuple36533USEDMULTIPLEtuple[1])), .store_ready(f1_store_ready), .load_ready_downstream(AO_ready), .load_ready(f1_load_ready), .load_reset(reset), .store_input(left_process_output), .store_output(f1_store_output));
  LiftHandshake_RunIffReady_LiftDecimate_fifo_SIZE128_uint8_Wnil_Hnil_Tnil_BYTES128 #(.INSTANCE_NAME({INSTANCE_NAME,"_f2"})) f2(.CLK(CLK), .load_input(unnamedtuple36395USEDMULTIPLEtuple), .load_output(f2_load_output), .store_reset(reset), .store_ready_downstream((unnamedtuple36533USEDMULTIPLEtuple[2])), .store_ready(f2_store_ready), .load_ready_downstream(AOr_ready), .load_ready(f2_load_ready), .load_reset(reset), .store_input(right_process_output), .store_output(f2_store_output));
  LiftHandshake_RunIffReady_LiftDecimate_fifo_SIZE128__uint8_uint16__Wnil_Hnil_Tnil_BYTES384 #(.INSTANCE_NAME({INSTANCE_NAME,"_f3"})) f3(.CLK(CLK), .load_input(unnamedtuple36395USEDMULTIPLEtuple), .load_output(f3_load_output), .store_reset(reset), .store_ready_downstream((unnamedtuple36533USEDMULTIPLEtuple[3])), .store_ready(f3_store_ready), .load_ready_downstream(display_ready), .load_ready(f3_load_ready), .load_reset(reset), .store_input(AM_process_output), .store_output(f3_store_output));
  MakeHandshake_displayOutput #(.INSTANCE_NAME({INSTANCE_NAME,"_display"})) display(.CLK(CLK), .ready_downstream(CRP_ready), .ready(display_ready), .reset(reset), .process_input(f3_load_output), .process_output(display_process_output));
  LiftHandshake_LiftDecimate_liftXYSeq_lift_CropSeq_uint8_4_1__W831_H495_T1 #(.INSTANCE_NAME({INSTANCE_NAME,"_CRP"})) CRP(.CLK(CLK), .ready_downstream(incrate_ready), .ready(CRP_ready), .reset(reset), .process_input(display_process_output), .process_output(CRP_process_output));
  LiftHandshake_WaitOnInput_ChangeRate_uint8_4_1__from1_to2_H1 #(.INSTANCE_NAME({INSTANCE_NAME,"_incrate"})) incrate(.CLK(CLK), .ready_downstream((unnamedtuple36533USEDMULTIPLEtuple[0])), .ready(incrate_ready), .reset(reset), .process_input(CRP_process_output), .process_output(incrate_process_output));
  LiftHandshake_WaitOnInput_ChangeRate_uint8_2_1__from4_to1_H1 #(.INSTANCE_NAME({INSTANCE_NAME,"_reducerate"})) reducerate(.CLK(CLK), .ready_downstream(pad_ready), .ready(reducerate_ready), .reset(reset), .process_input(process_input), .process_output(reducerate_process_output));
  LiftHandshake_WaitOnInput_PadSeq_uint8_2_1__W640_H480_L191_R0_B7_Top8_T11 #(.INSTANCE_NAME({INSTANCE_NAME,"_pad"})) pad(.CLK(CLK), .ready_downstream(oi0_ready), .ready(pad_ready), .reset(reset), .process_input(reducerate_process_output), .process_output(pad_process_output));
  MakeHandshake_slice_typeuint8_2_1__1_1__xl0_xh0_yl0_yh0 #(.INSTANCE_NAME({INSTANCE_NAME,"_oi0"})) oi0(.CLK(CLK), .ready_downstream(inp_broadcast_ready), .ready(oi0_ready), .reset(reset), .process_input(pad_process_output), .process_output(oi0_process_output));
  BroadcastStream_uint8_2_1__2 #(.INSTANCE_NAME({INSTANCE_NAME,"_inp_broadcast"})) inp_broadcast(.CLK(CLK), .ready_downstream({right_ready,left_ready}), .ready(inp_broadcast_ready), .reset_valid(reset), .process_input(oi0_process_output), .process_output(inp_broadcast_process_output));
  MakeHandshake_slice_typeuint8_2_1__xl0_xh0_yl0_yh0 #(.INSTANCE_NAME({INSTANCE_NAME,"_left"})) left(.CLK(CLK), .ready_downstream(f1_store_ready), .ready(left_ready), .reset(reset), .process_input(({inp_broadcast_process_output[16:0]})), .process_output(left_process_output));
  MakeHandshake_slice_typeuint8_2_1__xl1_xh1_yl0_yh0 #(.INSTANCE_NAME({INSTANCE_NAME,"_right"})) right(.CLK(CLK), .ready_downstream(f2_store_ready), .ready(right_ready), .reset(reset), .process_input(({inp_broadcast_process_output[33:17]})), .process_output(right_process_output));
  MakeHandshake_arrayop_uint8_W1_Hnil #(.INSTANCE_NAME({INSTANCE_NAME,"_AO"})) AO(.CLK(CLK), .ready_downstream(LB_ready), .ready(AO_ready), .reset(reset), .process_input(f1_load_output), .process_output(AO_process_output));
  stencilLinebufferPartialOverlap #(.INSTANCE_NAME({INSTANCE_NAME,"_LB"})) LB(.CLK(CLK), .ready_downstream(llb_ready), .ready(LB_ready), .reset(reset), .process_input(AO_process_output), .process_output(LB_process_output));
  MakeHandshake_unpackStencil_uint8_W16_H16_T2 #(.INSTANCE_NAME({INSTANCE_NAME,"_llb"})) llb(.CLK(CLK), .ready_downstream((merge_ready[0])), .ready(llb_ready), .reset(reset), .process_input(LB_process_output), .process_output(llb_process_output));
  MakeHandshake_arrayop_uint8_W1_Hnil #(.INSTANCE_NAME({INSTANCE_NAME,"_AOr"})) AOr(.CLK(CLK), .ready_downstream(rightLB_ready), .ready(AOr_ready), .reset(reset), .process_input(f2_load_output), .process_output(AOr_process_output));
  MakeHandshake_stencilLinebuffer_Auint8_w831_h495_xmin15_ymin15 #(.INSTANCE_NAME({INSTANCE_NAME,"_rightLB"})) rightLB(.CLK(CLK), .ready_downstream(rAO_ready), .ready(rightLB_ready), .reset(reset), .process_input(AOr_process_output), .process_output(rightLB_process_output));
  MakeHandshake_arrayop_uint8_16_16__W1_Hnil #(.INSTANCE_NAME({INSTANCE_NAME,"_rAO"})) rAO(.CLK(CLK), .ready_downstream(rup_ready), .ready(rAO_ready), .reset(reset), .process_input(rightLB_process_output), .process_output(rAO_process_output));
  LiftHandshake_WaitOnInput_UpsampleXSeq #(.INSTANCE_NAME({INSTANCE_NAME,"_rup"})) rup(.CLK(CLK), .ready_downstream(right2_ready), .ready(rup_ready), .reset(reset), .process_input(rAO_process_output), .process_output(rup_process_output));
  MakeHandshake_slice_typeuint8_16_16__1_1__xl0_xh0_yl0_yh0 #(.INSTANCE_NAME({INSTANCE_NAME,"_right2"})) right2(.CLK(CLK), .ready_downstream(rb2_ready), .ready(right2_ready), .reset(reset), .process_input(rup_process_output), .process_output(right2_process_output));
  MakeHandshake_Broadcast_2 #(.INSTANCE_NAME({INSTANCE_NAME,"_rb2"})) rb2(.CLK(CLK), .ready_downstream((merge_ready[1])), .ready(rb2_ready), .reset(reset), .process_input(right2_process_output), .process_output(rb2_process_output));
  SoAtoAoSHandshake_W2_H1_table__0x42b86538 #(.INSTANCE_NAME({INSTANCE_NAME,"_merge"})) merge(.CLK(CLK), .ready_downstream(mer_ready), .ready(merge_ready), .reset(reset), .process_input({rb2_process_output,llb_process_output}), .process_output(merge_process_output));
  MakeHandshake_map_packTupleArrays_table__0x4293c570_W2_H1 #(.INSTANCE_NAME({INSTANCE_NAME,"_mer"})) mer(.CLK(CLK), .ready_downstream(AM_ready), .ready(mer_ready), .reset(reset), .process_input(merge_process_output), .process_output(mer_process_output));
  LiftHandshake_LiftDecimate_argmin #(.INSTANCE_NAME({INSTANCE_NAME,"_AM"})) AM(.CLK(CLK), .ready_downstream(f3_store_ready), .ready(AM_ready), .reset(reset), .process_input(mer_process_output), .process_output(AM_process_output));
endmodule

module Overflow_153600(input CLK, input process_valid, input CE, input [63:0] process_input, output [64:0] process_output, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  reg [63:0] process_input_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin process_input_delay1_validunnamednull0_CECE <= process_input; end end
  wire [31:0] cnt_GET_OUTPUT;
  reg unnamedbinop36752_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedbinop36752_delay1_validunnamednull0_CECE <= {((cnt_GET_OUTPUT)<((32'd153600)))}; end end
  wire [31:0] cnt_SETBY_OUTPUT;
  assign process_output = {unnamedbinop36752_delay1_validunnamednull0_CECE,process_input_delay1_validunnamednull0_CECE};
  // function: process pure=false delay=1
  // function: reset pure=false delay=0
  RegBy_incif_1uint32_CEtable__0x45fd16f0_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_cnt"})) cnt(.CLK(CLK), .set_valid(reset), .CE(CE), .set_inp((32'd0)), .setby_valid(process_valid), .setby_inp((1'd1)), .SETBY_OUTPUT(cnt_SETBY_OUTPUT), .GET_OUTPUT(cnt_GET_OUTPUT));
endmodule

module LiftDecimate_Overflow_153600(input CLK, output ready, input reset, input CE, input process_valid, input [64:0] process_input, output [64:0] process_output);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(process_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'process'", INSTANCE_NAME);  end end
  assign ready = (1'd1);
  wire unnamedcast36780USEDMULTIPLEcast;assign unnamedcast36780USEDMULTIPLEcast = (process_input[64]); 
  wire [64:0] LiftDecimate_process_output;
  reg [63:0] unnamedcast36783_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast36783_delay1_validunnamednull0_CECE <= (LiftDecimate_process_output[63:0]); end end
  reg unnamedcast36780_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedcast36780_delay1_validunnamednull0_CECE <= unnamedcast36780USEDMULTIPLEcast; end end
  reg unnamedbinop36788_delay1_validunnamednull0_CECE;  always @ (posedge CLK) begin if (CE) begin unnamedbinop36788_delay1_validunnamednull0_CECE <= {((LiftDecimate_process_output[64])&&unnamedcast36780_delay1_validunnamednull0_CECE)}; end end
  assign process_output = {unnamedbinop36788_delay1_validunnamednull0_CECE,unnamedcast36783_delay1_validunnamednull0_CECE};
  // function: ready pure=true delay=0
  // function: reset pure=false delay=0
  // function: process pure=false delay=2
  Overflow_153600 #(.INSTANCE_NAME({INSTANCE_NAME,"_LiftDecimate"})) LiftDecimate(.CLK(CLK), .process_valid({(unnamedcast36780USEDMULTIPLEcast&&process_valid)}), .CE(CE), .process_input((process_input[63:0])), .process_output(LiftDecimate_process_output), .reset(reset));
endmodule

module ShiftRegister_2_CEtrue_TY1(input CLK, input pushPop_valid, input CE, input sr_input, output pushPop_out, input reset);
parameter INSTANCE_NAME="INST";
always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'pushPop'", INSTANCE_NAME);  end end
always @(posedge CLK) begin if(reset===1'bx) begin $display("Valid bit can't be x! Module '%s' function 'reset'", INSTANCE_NAME);  end end
  reg SR2;
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR1' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR1' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR1' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate36855USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate36855USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(sr_input):((1'd0)))}; 
  reg SR1;  always @ (posedge CLK) begin if ((unnamedcallArbitrate36855USEDMULTIPLEcallArbitrate[1]) && CE) begin SR1 <= (unnamedcallArbitrate36855USEDMULTIPLEcallArbitrate[0]); end end
  always @(posedge CLK) begin if(pushPop_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR2' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(reset===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'SR2' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,pushPop_valid})+({4'b0,reset})) > 5'd1) begin $display("error, function 'set' on instance 'SR2' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [1:0] unnamedcallArbitrate36861USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate36861USEDMULTIPLEcallArbitrate = {(pushPop_valid||reset),((pushPop_valid)?(SR1):((1'd0)))}; 
    always @ (posedge CLK) begin if ((unnamedcallArbitrate36861USEDMULTIPLEcallArbitrate[1]) && CE) begin SR2 <= (unnamedcallArbitrate36861USEDMULTIPLEcallArbitrate[0]); end end
  assign pushPop_out = SR2;
  // function: pushPop pure=false delay=0
  // function: reset pure=false delay=0
endmodule

module LiftHandshake_LiftDecimate_Overflow_153600(input CLK, input ready_downstream, output ready, input reset, input [64:0] process_input, output [64:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire inner_LiftDecimate_Overflow_153600_ready;
  assign ready = {(inner_LiftDecimate_Overflow_153600_ready&&ready_downstream)};
  wire unnamedbinop36825USEDMULTIPLEbinop;assign unnamedbinop36825USEDMULTIPLEbinop = {(reset||ready_downstream)}; 
  wire unnamedunary36826USEDMULTIPLEunary;assign unnamedunary36826USEDMULTIPLEunary = {(~reset)}; 
  wire [64:0] inner_LiftDecimate_Overflow_153600_process_output;
  wire validBitDelay_LiftDecimate_Overflow_153600_pushPop_out;
  wire [64:0] unnamedtuple36875USEDMULTIPLEtuple;assign unnamedtuple36875USEDMULTIPLEtuple = {{((inner_LiftDecimate_Overflow_153600_process_output[64])&&validBitDelay_LiftDecimate_Overflow_153600_pushPop_out)},(inner_LiftDecimate_Overflow_153600_process_output[63:0])}; 
  always @(posedge CLK) begin if({(~{((unnamedtuple36875USEDMULTIPLEtuple[64])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: output valid bit should not be X!",INSTANCE_NAME); end end
  always @(posedge CLK) begin if({(~{((process_input[64])===1'bx)})} == 1'b0 && (1'd1)==1'b1) begin $display("%s: LiftHandshake: input valid bit should not be X!",INSTANCE_NAME); end end
  assign process_output = unnamedtuple36875USEDMULTIPLEtuple;
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  LiftDecimate_Overflow_153600 #(.INSTANCE_NAME({INSTANCE_NAME,"_inner_LiftDecimate_Overflow_153600"})) inner_LiftDecimate_Overflow_153600(.CLK(CLK), .ready(inner_LiftDecimate_Overflow_153600_ready), .reset(reset), .CE(unnamedbinop36825USEDMULTIPLEbinop), .process_valid(unnamedunary36826USEDMULTIPLEunary), .process_input(process_input), .process_output(inner_LiftDecimate_Overflow_153600_process_output));
  ShiftRegister_2_CEtrue_TY1 #(.INSTANCE_NAME({INSTANCE_NAME,"_validBitDelay_LiftDecimate_Overflow_153600"})) validBitDelay_LiftDecimate_Overflow_153600(.CLK(CLK), .pushPop_valid(unnamedunary36826USEDMULTIPLEunary), .CE(unnamedbinop36825USEDMULTIPLEbinop), .sr_input((1'd1)), .pushPop_out(validBitDelay_LiftDecimate_Overflow_153600_pushPop_out), .reset(reset));
endmodule

module Underflow_Auint8_4_1__2_1__count153600_cycles6087906_toosoonnil_USfalse(input CLK, input ready_downstream, output ready, input reset, input [64:0] process_input, output [64:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  assign ready = ready_downstream;
  wire unnamedbinop37634USEDMULTIPLEbinop;assign unnamedbinop37634USEDMULTIPLEbinop = {(ready_downstream||reset)}; 
  wire [31:0] cycleCount_GET_OUTPUT;
  wire unnamedbinop37633USEDMULTIPLEbinop;assign unnamedbinop37633USEDMULTIPLEbinop = {((cycleCount_GET_OUTPUT)>((32'd6087906)))}; 
  wire [31:0] outputCount_GET_OUTPUT;
  wire unnamedcast37627USEDMULTIPLEcast;assign unnamedcast37627USEDMULTIPLEcast = (process_input[64]); 
  wire unnamedunary37653USEDMULTIPLEunary;assign unnamedunary37653USEDMULTIPLEunary = {(~reset)}; 
  wire [31:0] outputCount_SETBY_OUTPUT;
  wire [31:0] cycleCount_SETBY_OUTPUT;
  assign process_output = {{({({(unnamedbinop37633USEDMULTIPLEbinop&&{((outputCount_GET_OUTPUT)<((32'd153600)))})}||{({(~unnamedbinop37633USEDMULTIPLEbinop)}&&unnamedcast37627USEDMULTIPLEcast)})}&&unnamedunary37653USEDMULTIPLEunary)},((unnamedbinop37633USEDMULTIPLEbinop)?((64'd3735928559)):((process_input[63:0])))};
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  RegBy_incif_1uint32_CEtable__0x45fd16f0_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_outputCount"})) outputCount(.CLK(CLK), .set_valid(reset), .CE(unnamedbinop37634USEDMULTIPLEbinop), .set_inp((32'd0)), .setby_valid(unnamedunary37653USEDMULTIPLEunary), .setby_inp({(ready_downstream&&{(unnamedcast37627USEDMULTIPLEcast||unnamedbinop37633USEDMULTIPLEbinop)})}), .SETBY_OUTPUT(outputCount_SETBY_OUTPUT), .GET_OUTPUT(outputCount_GET_OUTPUT));
  RegBy_incif_1uint32_CEtable__0x45fd16f0_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_cycleCount"})) cycleCount(.CLK(CLK), .set_valid(reset), .CE(unnamedbinop37634USEDMULTIPLEbinop), .set_inp((32'd0)), .setby_valid(unnamedunary37653USEDMULTIPLEunary), .setby_inp((1'd1)), .SETBY_OUTPUT(cycleCount_SETBY_OUTPUT), .GET_OUTPUT(cycleCount_GET_OUTPUT));
endmodule

module incif_wrapuint32_153615_inc1(input CLK, input CE, input [32:0] process_input, output [31:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [31:0] unnamedcast37311USEDMULTIPLEcast;assign unnamedcast37311USEDMULTIPLEcast = (process_input[31:0]); 
  assign process_output = (((process_input[32]))?((({(unnamedcast37311USEDMULTIPLEcast==(32'd153615))})?((32'd0)):({(unnamedcast37311USEDMULTIPLEcast+(32'd1))}))):(unnamedcast37311USEDMULTIPLEcast));
  // function: process pure=true delay=0
endmodule

module RegBy_incif_wrapuint32_153615_inc1_CEtrue_initnil(input CLK, input set_valid, input CE, input [31:0] set_inp, input setby_valid, input setby_inp, output [31:0] SETBY_OUTPUT, output [31:0] GET_OUTPUT);
parameter INSTANCE_NAME="INST";
  reg [31:0] R;
  wire [31:0] regby_inner_process_output;
  always @(posedge CLK) begin if(set_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(setby_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,set_valid})+({4'b0,setby_valid})) > 5'd1) begin $display("error, function 'set' on instance 'R' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [32:0] unnamedcallArbitrate37362USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate37362USEDMULTIPLEcallArbitrate = {(set_valid||setby_valid),((set_valid)?(set_inp):(regby_inner_process_output))}; 
    always @ (posedge CLK) begin if ((unnamedcallArbitrate37362USEDMULTIPLEcallArbitrate[32]) && CE) begin R <= (unnamedcallArbitrate37362USEDMULTIPLEcallArbitrate[31:0]); end end
  assign SETBY_OUTPUT = regby_inner_process_output;
  assign GET_OUTPUT = R;
  // function: set pure=false ONLY WIRE
  // function: setby pure=false ONLY WIRE
  // function: get pure=true ONLY WIRE
  incif_wrapuint32_153615_inc1 #(.INSTANCE_NAME({INSTANCE_NAME,"_regby_inner"})) regby_inner(.CLK(CLK), .CE(CE), .process_input({setby_inp,R}), .process_output(regby_inner_process_output));
endmodule

module incif_1uint32_CEnil(input CLK, input [32:0] process_input, output [31:0] process_output);
parameter INSTANCE_NAME="INST";
  wire [31:0] unnamedcast37371USEDMULTIPLEcast;assign unnamedcast37371USEDMULTIPLEcast = (process_input[31:0]); 
  assign process_output = (((process_input[32]))?({(unnamedcast37371USEDMULTIPLEcast+(32'd1))}):(unnamedcast37371USEDMULTIPLEcast));
  // function: process pure=true delay=0
endmodule

module RegBy_incif_1uint32_CEnil_CEfalse_initnil(input CLK, input set_valid, input [31:0] set_inp, input setby_valid, input setby_inp, output [31:0] SETBY_OUTPUT, output [31:0] GET_OUTPUT);
parameter INSTANCE_NAME="INST";
  reg [31:0] R;
  wire [31:0] regby_inner_process_output;
  always @(posedge CLK) begin if(set_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if(setby_valid===1'bx) begin $display("valid bit can't be x! Module '%s' instance 'R' function 'set'", INSTANCE_NAME); end end
  always @(posedge CLK) begin if((({4'b0,set_valid})+({4'b0,setby_valid})) > 5'd1) begin $display("error, function 'set' on instance 'R' in module '%s' has multiple valid bits active in same cycle!",INSTANCE_NAME);$finish(); end end
  wire [32:0] unnamedcallArbitrate37403USEDMULTIPLEcallArbitrate;assign unnamedcallArbitrate37403USEDMULTIPLEcallArbitrate = {(set_valid||setby_valid),((set_valid)?(set_inp):(regby_inner_process_output))}; 
    always @ (posedge CLK) begin R <= (unnamedcallArbitrate37403USEDMULTIPLEcallArbitrate[31:0]); end
  assign SETBY_OUTPUT = regby_inner_process_output;
  assign GET_OUTPUT = R;
  // function: set pure=false ONLY WIRE
  // function: setby pure=false ONLY WIRE
  // function: get pure=true ONLY WIRE
  incif_1uint32_CEnil #(.INSTANCE_NAME({INSTANCE_NAME,"_regby_inner"})) regby_inner(.CLK(CLK), .process_input({setby_inp,R}), .process_output(regby_inner_process_output));
endmodule

module CycleCounter_Auint8_4_1__2_1__count153600(input CLK, input ready_downstream, output ready, input reset, input [64:0] process_input, output [64:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire [31:0] outputCount_GET_OUTPUT;
  wire unnamedbinop37416USEDMULTIPLEbinop;assign unnamedbinop37416USEDMULTIPLEbinop = {((outputCount_GET_OUTPUT)>=((32'd153600)))}; 
  wire unnamedunary37439USEDMULTIPLEunary;assign unnamedunary37439USEDMULTIPLEunary = {(~unnamedbinop37416USEDMULTIPLEbinop)}; 
  assign ready = {(ready_downstream&&unnamedunary37439USEDMULTIPLEunary)};
  wire unnamedbinop37417USEDMULTIPLEbinop;assign unnamedbinop37417USEDMULTIPLEbinop = {(ready_downstream||reset)}; 
  wire [31:0] cycleCount_GET_OUTPUT;
  wire unnamedcast37410USEDMULTIPLEcast;assign unnamedcast37410USEDMULTIPLEcast = (process_input[64]); 
  wire unnamedunary37432USEDMULTIPLEunary;assign unnamedunary37432USEDMULTIPLEunary = {(~reset)}; 
  wire [31:0] outputCount_SETBY_OUTPUT;
  wire [31:0] cycleCount_SETBY_OUTPUT;
  assign process_output = {{({(unnamedbinop37416USEDMULTIPLEbinop||unnamedcast37410USEDMULTIPLEcast)}&&unnamedunary37432USEDMULTIPLEunary)},((unnamedbinop37416USEDMULTIPLEbinop)?({cycleCount_GET_OUTPUT,cycleCount_GET_OUTPUT}):((process_input[63:0])))};
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  RegBy_incif_wrapuint32_153615_inc1_CEtrue_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_outputCount"})) outputCount(.CLK(CLK), .set_valid(reset), .CE(unnamedbinop37417USEDMULTIPLEbinop), .set_inp((32'd0)), .setby_valid(unnamedunary37432USEDMULTIPLEunary), .setby_inp({(ready_downstream&&{(unnamedcast37410USEDMULTIPLEcast||unnamedbinop37416USEDMULTIPLEbinop)})}), .SETBY_OUTPUT(outputCount_SETBY_OUTPUT), .GET_OUTPUT(outputCount_GET_OUTPUT));
  RegBy_incif_1uint32_CEnil_CEfalse_initnil #(.INSTANCE_NAME({INSTANCE_NAME,"_cycleCount"})) cycleCount(.CLK(CLK), .set_valid(reset), .set_inp((32'd0)), .setby_valid(unnamedunary37432USEDMULTIPLEunary), .setby_inp(unnamedunary37439USEDMULTIPLEunary), .SETBY_OUTPUT(cycleCount_SETBY_OUTPUT), .GET_OUTPUT(cycleCount_GET_OUTPUT));
endmodule

module harnessaxi(input CLK, input ready_downstream, output ready, input reset, input [64:0] process_input, output [64:0] process_output);
parameter INSTANCE_NAME="INST";
parameter OUTPUT_COUNT=0;
parameter INPUT_COUNT=0;
  wire cycleCounter_ready;
  wire underflow_ready;
  wire overflow_ready;
  wire hsfna_ready;
  wire underflow_US_ready;
  assign ready = underflow_US_ready;
  wire [64:0] underflow_US_process_output;
  wire [64:0] hsfna_process_output;
  wire [64:0] overflow_process_output;
  wire [64:0] underflow_process_output;
  wire [64:0] cycleCounter_process_output;
  assign process_output = cycleCounter_process_output;
  // function: ready pure=true ONLY WIRE
  // function: reset pure=false ONLY WIRE
  // function: process pure=false ONLY WIRE
  Underflow_Auint8_2_1__4_1__count76800_cycles6087906_toosoonnil_UStrue #(.INSTANCE_NAME({INSTANCE_NAME,"_underflow_US"})) underflow_US(.CLK(CLK), .ready_downstream(hsfna_ready), .ready(underflow_US_ready), .reset(reset), .process_input(process_input), .process_output(underflow_US_process_output));
  hsfn #(.INSTANCE_NAME({INSTANCE_NAME,"_hsfna"})) hsfna(.CLK(CLK), .ready_downstream(overflow_ready), .ready(hsfna_ready), .reset(reset), .process_input(underflow_US_process_output), .process_output(hsfna_process_output));
  LiftHandshake_LiftDecimate_Overflow_153600 #(.INSTANCE_NAME({INSTANCE_NAME,"_overflow"})) overflow(.CLK(CLK), .ready_downstream(underflow_ready), .ready(overflow_ready), .reset(reset), .process_input(hsfna_process_output), .process_output(overflow_process_output));
  Underflow_Auint8_4_1__2_1__count153600_cycles6087906_toosoonnil_USfalse #(.INSTANCE_NAME({INSTANCE_NAME,"_underflow"})) underflow(.CLK(CLK), .ready_downstream(cycleCounter_ready), .ready(underflow_ready), .reset(reset), .process_input(overflow_process_output), .process_output(underflow_process_output));
  CycleCounter_Auint8_4_1__2_1__count153600 #(.INSTANCE_NAME({INSTANCE_NAME,"_cycleCounter"})) cycleCounter(.CLK(CLK), .ready_downstream(ready_downstream), .ready(cycleCounter_ready), .reset(reset), .process_input(underflow_process_output), .process_output(cycleCounter_process_output));
endmodule

`timescale 1ps/1ps

module ict106_axilite_conv2 #
  (
   parameter integer C_AXI_ID_WIDTH              = 12,
   parameter integer C_AXI_ADDR_WIDTH            = 32,
   parameter integer C_AXI_DATA_WIDTH            = 32 // CONSTANT
   )
  (
   // System Signals
   input  wire                          ACLK,
   input  wire                          ARESETN,
   input  wire [C_AXI_ID_WIDTH-1:0]     S_AXI_AWID,
   input  wire [C_AXI_ADDR_WIDTH-1:0]   S_AXI_AWADDR,
   input  wire                          S_AXI_AWVALID,
   output wire                          S_AXI_AWREADY,
   input  wire [C_AXI_DATA_WIDTH-1:0]   S_AXI_WDATA,
   input  wire [C_AXI_DATA_WIDTH/8-1:0] S_AXI_WSTRB,
   input  wire                          S_AXI_WVALID,
   output wire                          S_AXI_WREADY,
   output wire [C_AXI_ID_WIDTH-1:0]     S_AXI_BID,
   output wire [2-1:0]                  S_AXI_BRESP,
   output wire                          S_AXI_BVALID,
   input  wire                          S_AXI_BREADY,
   input  wire [C_AXI_ID_WIDTH-1:0]     S_AXI_ARID,
   input  wire [C_AXI_ADDR_WIDTH-1:0]   S_AXI_ARADDR,
   input  wire                          S_AXI_ARVALID,
   output wire                          S_AXI_ARREADY,
   output wire [C_AXI_ID_WIDTH-1:0]     S_AXI_RID,
   output wire [C_AXI_DATA_WIDTH-1:0]   S_AXI_RDATA,
   output wire [2-1:0]                  S_AXI_RRESP,
   output wire                          S_AXI_RLAST,    // Constant =1
   output wire                          S_AXI_RVALID,
   input  wire                          S_AXI_RREADY,
   output wire [C_AXI_ADDR_WIDTH-1:0]   M_AXI_AWADDR,
   output wire                          M_AXI_AWVALID,
   input  wire                          M_AXI_AWREADY,
   output wire [C_AXI_DATA_WIDTH-1:0]   M_AXI_WDATA,
   output wire [C_AXI_DATA_WIDTH/8-1:0] M_AXI_WSTRB,
   output wire                          M_AXI_WVALID,
   input  wire                          M_AXI_WREADY,
   input  wire [2-1:0]                  M_AXI_BRESP,
   input  wire                          M_AXI_BVALID,
   output wire                          M_AXI_BREADY,
   output wire [C_AXI_ADDR_WIDTH-1:0]   M_AXI_ARADDR,
   output wire                          M_AXI_ARVALID,
   input  wire                          M_AXI_ARREADY,
   input  wire [C_AXI_DATA_WIDTH-1:0]   M_AXI_RDATA,
   input  wire [2-1:0]                  M_AXI_RRESP,
   input  wire                          M_AXI_RVALID,
   output wire                          M_AXI_RREADY
  );
  
  wire [31:0] m_axaddr;

  // Arbiter
  reg read_active;
  reg write_active;
  reg busy;

  wire read_req;
  wire write_req;
  wire read_complete;
  wire write_complete;
  
  reg [1:0] areset_d; // Reset delay register
  always @(posedge ACLK) begin
    areset_d <= {areset_d[0], ~ARESETN};
  end
  
  assign read_req  = S_AXI_ARVALID & ~write_active & ~busy & ~|areset_d;
  assign write_req = (S_AXI_AWVALID & ~read_active & ~busy & ~S_AXI_ARVALID & ~|areset_d) | (write_active & ~busy);

  assign read_complete  = M_AXI_RVALID & S_AXI_RREADY;
  assign write_complete = M_AXI_BVALID & S_AXI_BREADY;

  always @(posedge ACLK) begin : arbiter_read_ff
    if (~ARESETN)
      read_active <= 1'b0;
    else if (read_complete)
      read_active <= 1'b0;
    else if (read_req)
      read_active <= 1'b1;
  end

  always @(posedge ACLK) begin : arbiter_write_ff
    if (~ARESETN)
      write_active <= 1'b0;
    else if (write_complete)
      write_active <= 1'b0;
    else if (write_req)
      write_active <= 1'b1;
  end

  always @(posedge ACLK) begin : arbiter_busy_ff
    if (~ARESETN)
      busy <= 1'b0;
    else if (read_complete | write_complete)
      busy <= 1'b0;
    else if ((S_AXI_AWVALID & M_AXI_AWREADY & ~read_req) | (S_AXI_ARVALID & M_AXI_ARREADY & ~write_req))
      busy <= 1'b1;
  end

  assign M_AXI_ARVALID = read_req;
  assign S_AXI_ARREADY = M_AXI_ARREADY & read_req;

  assign M_AXI_AWVALID = write_req;
  assign S_AXI_AWREADY = M_AXI_AWREADY & write_req;

  assign M_AXI_RREADY  = S_AXI_RREADY & read_active;
  assign S_AXI_RVALID  = M_AXI_RVALID & read_active;

  assign M_AXI_BREADY  = S_AXI_BREADY & write_active;
  assign S_AXI_BVALID  = M_AXI_BVALID & write_active;

  // Address multiplexer
  assign m_axaddr = (read_req) ? S_AXI_ARADDR : S_AXI_AWADDR;

  // Id multiplexer and flip-flop
  reg [C_AXI_ID_WIDTH-1:0] s_axid;

  always @(posedge ACLK) begin : axid
    if      (~ARESETN)    s_axid <= {C_AXI_ID_WIDTH{1'b0}};
    else if (read_req)  s_axid <= S_AXI_ARID;
    else if (write_req) s_axid <= S_AXI_AWID;
  end

  assign S_AXI_BID = s_axid;
  assign S_AXI_RID = s_axid;

  assign M_AXI_AWADDR = m_axaddr;
  assign M_AXI_ARADDR = m_axaddr;


  // Feed-through signals
  assign S_AXI_WREADY   = M_AXI_WREADY & ~|areset_d;
  assign S_AXI_BRESP    = M_AXI_BRESP;
  assign S_AXI_RDATA    = M_AXI_RDATA;
  assign S_AXI_RRESP    = M_AXI_RRESP;
  assign S_AXI_RLAST    = 1'b1;

  assign M_AXI_WVALID   = S_AXI_WVALID & ~|areset_d;
  assign M_AXI_WDATA    = S_AXI_WDATA;
  assign M_AXI_WSTRB    = S_AXI_WSTRB;

endmodule

module Conf(
    input ACLK,
    input ARESETN,
    //AXI Inputs
    input [31:0] S_AXI_ARADDR,
    input [11:0] S_AXI_ARID,
    output S_AXI_ARREADY,
    input S_AXI_ARVALID,
    input [31:0] S_AXI_AWADDR,
    input [11:0] S_AXI_AWID,
    output S_AXI_AWREADY,
    input S_AXI_AWVALID,
    output [11:0] S_AXI_BID,
    input S_AXI_BREADY,
    output [1:0] S_AXI_BRESP,
    output S_AXI_BVALID,
    output [31:0] S_AXI_RDATA,
    output [11:0] S_AXI_RID,
    output S_AXI_RLAST,
    input S_AXI_RREADY,
    output [1:0] S_AXI_RRESP,
    output S_AXI_RVALID,
    input [31:0] S_AXI_WDATA,
    output S_AXI_WREADY,
    input [3:0] S_AXI_WSTRB,
    input S_AXI_WVALID,
    
    output CONFIG_VALID,
    input CONFIG_READY,
    output [31:0] CONFIG_CMD,
    output [31:0] CONFIG_SRC,
    output [31:0] CONFIG_DEST,
    output [31:0] CONFIG_LEN,
    output CONFIG_IRQ
    );

    //Convert Input signals to AXI lite, to avoid ID matching
    wire [31:0] LITE_ARADDR;
    wire LITE_ARREADY;
    wire LITE_ARVALID;
    wire [31:0] LITE_AWADDR;
    wire LITE_AWREADY;
    wire LITE_AWVALID;
    wire LITE_BREADY;
    reg [1:0] LITE_BRESP;
    wire LITE_BVALID;
    reg [31:0] LITE_RDATA;
    wire LITE_RREADY;
    reg [1:0] LITE_RRESP;
    wire LITE_RVALID;
    wire [31:0] LITE_WDATA;
    wire LITE_WREADY;
    wire [3:0] LITE_WSTRB;
    wire LITE_WVALID;
    
    ict106_axilite_conv axilite(
    .ACLK(ACLK),
    .ARESETN(ARESETN),
    .S_AXI_ARADDR(S_AXI_ARADDR), 
    .S_AXI_ARID(S_AXI_ARID),  
    .S_AXI_ARREADY(S_AXI_ARREADY), 
    .S_AXI_ARVALID(S_AXI_ARVALID), 
    .S_AXI_AWADDR(S_AXI_AWADDR), 
    .S_AXI_AWID(S_AXI_AWID), 
    .S_AXI_AWREADY(S_AXI_AWREADY), 
    .S_AXI_AWVALID(S_AXI_AWVALID), 
    .S_AXI_BID(S_AXI_BID), 
    .S_AXI_BREADY(S_AXI_BREADY), 
    .S_AXI_BRESP(S_AXI_BRESP), 
    .S_AXI_BVALID(S_AXI_BVALID), 
    .S_AXI_RDATA(S_AXI_RDATA), 
    .S_AXI_RID(S_AXI_RID), 
    .S_AXI_RLAST(S_AXI_RLAST), 
    .S_AXI_RREADY(S_AXI_RREADY), 
    .S_AXI_RRESP(S_AXI_RRESP), 
    .S_AXI_RVALID(S_AXI_RVALID), 
    .S_AXI_WDATA(S_AXI_WDATA), 
    .S_AXI_WREADY(S_AXI_WREADY), 
    .S_AXI_WSTRB(S_AXI_WSTRB), 
    .S_AXI_WVALID(S_AXI_WVALID),
       
    .M_AXI_ARADDR(LITE_ARADDR),
    .M_AXI_ARREADY(LITE_ARREADY),
    .M_AXI_ARVALID(LITE_ARVALID),
    .M_AXI_AWADDR(LITE_AWADDR),
    .M_AXI_AWREADY(LITE_AWREADY),
    .M_AXI_AWVALID(LITE_AWVALID),
    .M_AXI_BREADY(LITE_BREADY),
    .M_AXI_BRESP(LITE_BRESP),
    .M_AXI_BVALID(LITE_BVALID),
    .M_AXI_RDATA(LITE_RDATA),
    .M_AXI_RREADY(LITE_RREADY),
    .M_AXI_RRESP(LITE_RRESP),
    .M_AXI_RVALID(LITE_RVALID),
    .M_AXI_WDATA(LITE_WDATA),
    .M_AXI_WREADY(LITE_WREADY),
    .M_AXI_WSTRB(LITE_WSTRB),
    .M_AXI_WVALID(LITE_WVALID)
  );

parameter NREG = 4;
parameter W = 32;

reg [W-1:0] data[NREG-1:0];

parameter IDLE = 0, RWAIT = 1;
parameter OK = 2'b00, SLVERR = 2'b10;

reg [31:0] counter;

//READS
reg r_state;
wire [1:0] r_select;
assign r_select  = LITE_ARADDR[3:2];
assign ar_good = {LITE_ARADDR[31:4], 2'b00, LITE_ARADDR[1:0]} == 32'h70000000;
assign LITE_ARREADY = (r_state == IDLE);
assign LITE_RVALID = (r_state == RWAIT);
always @(posedge ACLK) begin
    if(ARESETN == 0) begin
        r_state <= IDLE;
    end else case(r_state)
        IDLE: begin
            if(LITE_ARVALID) begin
                LITE_RRESP <= ar_good ? OK : SLVERR;
                LITE_RDATA <= (r_select == 2'b0) ? counter : data[r_select];
                r_state <= RWAIT;
            end
        end
        RWAIT: begin
            if(LITE_RREADY)
                r_state <= IDLE;
        end
    endcase
end 

//WRITES
reg w_state;
reg [1:0] w_select_r;
reg w_wrotedata;
reg w_wroteresp;

wire [1:0] w_select;
assign w_select  = LITE_AWADDR[3:2];
assign aw_good = {LITE_AWADDR[31:4], 2'b00, LITE_AWADDR[1:0]} == 32'h70000000;

assign LITE_AWREADY = (w_state == IDLE);
assign LITE_WREADY = (w_state == RWAIT) && !w_wrotedata;
assign LITE_BVALID = (w_state == RWAIT) && !w_wroteresp;

always @(posedge ACLK) begin
    if(ARESETN == 0) begin
        w_state <= IDLE;
        w_wrotedata <= 0;
        w_wroteresp <= 0;
    end else case(w_state)
        IDLE: begin
            if(LITE_AWVALID) begin
                LITE_BRESP <= aw_good ? OK : SLVERR;
                w_select_r <= w_select;
                w_state <= RWAIT; 
                w_wrotedata <= 0;
                w_wroteresp <= 0;
            end
        end
        RWAIT: begin
            if (LITE_WREADY)
                data[w_select_r] <= LITE_WDATA;
            if((w_wrotedata || LITE_WVALID) && (w_wroteresp || LITE_BREADY)) begin
                w_wrotedata <= 0;
                w_wroteresp <= 0;
                w_state <= IDLE;
            end else if (LITE_WVALID)
                w_wrotedata <= 1;
            else if (LITE_BREADY)
                w_wroteresp <= 1;
        end
    endcase
end

reg v_state;
assign CONFIG_VALID = (v_state == RWAIT);
always @(posedge ACLK) begin
    if (ARESETN == 0)
        v_state <= IDLE;
    else case(v_state)
        IDLE:
            if (LITE_WVALID && LITE_WREADY && w_select_r == 2'b00)
                v_state <= RWAIT;
        RWAIT:
            if (CONFIG_READY)
                v_state <= IDLE;
    endcase
end

assign CONFIG_CMD = data[0];
assign CONFIG_SRC = data[1];
assign CONFIG_DEST = data[2];
assign CONFIG_LEN = data[3];


//how many cycles does the operation take?
always @(posedge ACLK) begin
    if (ARESETN == 0)
        counter <= 0;
    else if (CONFIG_READY && CONFIG_VALID)
        counter <= 0;
    else if (!CONFIG_READY)
        counter <= counter + 1;
end

reg busy;
reg busy_last;
always @(posedge ACLK) begin
    if (ARESETN == 0) begin
        busy <= 0;
        busy_last <= 0;
    end else begin
        if (CONFIG_READY) begin
            busy <= CONFIG_VALID ? 1 : 0;
        end
        busy_last <= busy;
    end
end

assign CONFIG_IRQ = !busy;

endmodule // Conf

module DRAMReader(
    //AXI port
    input ACLK,
    input ARESETN,
    output reg [31:0] M_AXI_ARADDR,
    input M_AXI_ARREADY,
    output  M_AXI_ARVALID,
    input [63:0] M_AXI_RDATA,
    output M_AXI_RREADY,
    input [1:0] M_AXI_RRESP,
    input M_AXI_RVALID,
    input M_AXI_RLAST,
    output [3:0] M_AXI_ARLEN,
    output [1:0] M_AXI_ARSIZE,
    output [1:0] M_AXI_ARBURST,
    
    //Control config
    input CONFIG_VALID,
    output CONFIG_READY,
    input [31:0] CONFIG_START_ADDR,
    input [31:0] CONFIG_NBYTES,
    
    //RAM port
    input DATA_READY_DOWNSTREAM,
    output DATA_VALID,
    output [63:0] DATA
);

assign M_AXI_ARLEN = 4'b1111;
assign M_AXI_ARSIZE = 2'b11;
assign M_AXI_ARBURST = 2'b01;
parameter IDLE = 0, RWAIT = 1;
    
//ADDR logic
reg [31:0] a_count;
reg a_state;  
assign M_AXI_ARVALID = (a_state == RWAIT);
always @(posedge ACLK) begin
    if (ARESETN == 0) begin
        a_state <= IDLE;
        M_AXI_ARADDR <= 0;
        a_count <= 0;
    end else case(a_state)
        IDLE: begin
            if(CONFIG_VALID) begin
                M_AXI_ARADDR <= CONFIG_START_ADDR;
                a_count <= CONFIG_NBYTES[31:7];
                a_state <= RWAIT;
            end
        end
        RWAIT: begin
            if (M_AXI_ARREADY == 1) begin
                if(a_count - 1 == 0)
                    a_state <= IDLE;
                a_count <= a_count - 1;
                M_AXI_ARADDR <= M_AXI_ARADDR + 128; // Bursts are 128 bytes long
            end
        end
    endcase
end
    
//READ logic
reg [31:0] b_count;
reg r_state;
assign M_AXI_RREADY = (r_state == RWAIT) && DATA_READY_DOWNSTREAM;
always @(posedge ACLK) begin
    if (ARESETN == 0) begin
        r_state <= IDLE;
        b_count <= 0;
    end else case(r_state)
        IDLE: begin
            if(CONFIG_VALID) begin
                b_count <= {CONFIG_NBYTES[31:7],7'b0}; // round to nearest 128 bytes
                r_state <= RWAIT;
            end
        end
        RWAIT: begin
            if (M_AXI_RVALID && DATA_READY_DOWNSTREAM) begin
                //use M_AXI_RDATA
                if(b_count - 8 == 0)
                    r_state <= IDLE;
                b_count <= b_count - 8; // each valid cycle the bus provides 8 bytes
            end
        end
    endcase
end

assign DATA = M_AXI_RDATA;
assign DATA_VALID = M_AXI_RVALID && (r_state == RWAIT);
assign CONFIG_READY = (r_state == IDLE) && (a_state == IDLE);

endmodule // DRAMReader

module DRAMWriter(
    //AXI port
    input ACLK,
    input ARESETN,
    output reg [31:0] M_AXI_AWADDR,
    input M_AXI_AWREADY,
    output M_AXI_AWVALID,
    
    output [63:0] M_AXI_WDATA,
    output [7:0] M_AXI_WSTRB,
    input M_AXI_WREADY,
    output M_AXI_WVALID,
    output M_AXI_WLAST,
    
    input [1:0] M_AXI_BRESP,
    input M_AXI_BVALID,
    output M_AXI_BREADY,
    
    output [3:0] M_AXI_AWLEN,
    output [1:0] M_AXI_AWSIZE,
    output [1:0] M_AXI_AWBURST,
    
    //Control config
    input CONFIG_VALID,
    output CONFIG_READY,
    input [31:0] CONFIG_START_ADDR,
    input [31:0] CONFIG_NBYTES,
    
    //RAM port
    input [63:0] DATA,
    output DATA_READY,
    input DATA_VALID

);

assign M_AXI_AWLEN = 4'b1111;
assign M_AXI_AWSIZE = 2'b11;
assign M_AXI_AWBURST = 2'b01;
assign M_AXI_WSTRB = 8'b11111111;

parameter IDLE = 0, RWAIT = 1;
    
//ADDR logic
reg [31:0] a_count;
reg a_state;  
assign M_AXI_AWVALID = (a_state == RWAIT);
always @(posedge ACLK) begin
    if (ARESETN == 0) begin
        a_state <= IDLE;
        M_AXI_AWADDR <= 0;
        a_count <= 0;
    end else case(a_state)
        IDLE: begin
            if(CONFIG_VALID) begin
                M_AXI_AWADDR <= CONFIG_START_ADDR;
                a_count <= CONFIG_NBYTES[31:7];
                a_state <= RWAIT;
            end
        end
        RWAIT: begin
            if (M_AXI_AWREADY == 1) begin
                if(a_count - 1 == 0)
                    a_state <= IDLE;
                a_count <= a_count - 1;
                M_AXI_AWADDR <= M_AXI_AWADDR + 128; 
            end
        end
    endcase
end

//WRITE logic
reg [31:0] b_count;
reg w_state;
always @(posedge ACLK) begin
    if (ARESETN == 0) begin
        w_state <= IDLE;
        b_count <= 0;
    end else case(w_state)
        IDLE: begin
            if(CONFIG_VALID) begin
                b_count <= {CONFIG_NBYTES[31:7],7'b0};
                w_state <= RWAIT;
                last_count <= 4'b1111;
            end
        end
        RWAIT: begin
            if (M_AXI_WREADY && M_AXI_WVALID) begin
                //use M_AXI_WDATA
                if(b_count - 8 == 0) begin
                    w_state <= IDLE;
                end
                last_count <= last_count - 4'b1;
                b_count <= b_count - 8;
            end
        end
    endcase
end

reg [3:0] last_count;
assign M_AXI_WLAST = last_count == 4'b0000;

assign M_AXI_WVALID = (w_state == RWAIT) && DATA_VALID;

assign DATA_READY = (w_state == RWAIT) && M_AXI_WREADY;
   
assign CONFIG_READY = (w_state == IDLE) && (a_state == IDLE);

assign M_AXI_BREADY = 1;

assign M_AXI_WDATA = DATA;

endmodule // DRAMWriter

//-----------------------------------------------------------------------------
// system.v
//-----------------------------------------------------------------------------

// The axi bus expects the number of valid data items to exactly match the # of addresses we send.
// This module checks for underflow (too few valid data items). If there are too few, it inserts DEADBEEFs to make it correct.
// lengthOutput is in bytes
module UnderflowShim(input CLK, input RST, input [31:0] lengthOutput, input [63:0] inp, input inp_valid, output [63:0] out, output out_valid);
   parameter WAIT_CYCLES = 2048;
   
   reg [31:0] outCnt;
   reg [31:0] outLen;

   reg        fixupMode;
   reg [31:0]  outClks = 0;
   
   
   always@(posedge CLK) begin
     if (RST) begin 
        outCnt <= 32'd0;
        outLen <= lengthOutput;
        fixupMode <= 1'b0;
        outClks <= 32'd0;
     end else begin
        outClks <= outClks + 32'd1;
        
        if(inp_valid || fixupMode) begin outCnt <= outCnt+32'd8; end // AXI does 8 bytes per clock
        if(outClks > WAIT_CYCLES) begin fixupMode <= 1'b1; end
     end
   end

   assign out = (fixupMode)?(64'hDEAD):(inp);
   assign out_valid = (RST)?(1'b0):((fixupMode)?(outCnt<outLen):(inp_valid));
endmodule

module stage
  (
    inout [53:0] MIO,
    inout PS_SRSTB,
    inout PS_CLK,
    inout PS_PORB,
    inout DDR_Clk,
    inout DDR_Clk_n,
    inout DDR_CKE,
    inout DDR_CS_n,
    inout DDR_RAS_n,
    inout DDR_CAS_n,
    output DDR_WEB,
    inout [2:0] DDR_BankAddr,
    inout [14:0] DDR_Addr,
    inout DDR_ODT,
    inout DDR_DRSTB,
    inout [31:0] DDR_DQ,
    inout [3:0] DDR_DM,
    inout [3:0] DDR_DQS,
    inout [3:0] DDR_DQS_n,
    inout DDR_VRN,
    inout DDR_VRP,
    output [7:0] LED
  );

  wire [3:0] fclk;
  wire [3:0] fclkresetn;
  wire FCLK0;
  BUFG bufg(.I(fclk[0]),.O(FCLK0));
  assign ARESETN = fclkresetn[0];
  
  
    wire [31:0] PS7_ARADDR;
    wire [11:0] PS7_ARID;
    wire [2:0] PS7_ARPROT;
    wire PS7_ARREADY;
    wire PS7_ARVALID;
    wire [31:0] PS7_AWADDR;
    wire [11:0] PS7_AWID;
    wire [2:0] PS7_AWPROT;
    wire PS7_AWREADY;
    wire PS7_AWVALID;
    wire [11:0] PS7_BID;
    wire PS7_BREADY;
    wire [1:0] PS7_BRESP;
    wire PS7_BVALID;
    wire [31:0] PS7_RDATA;
    wire [11:0] PS7_RID;
    wire PS7_RLAST;
    wire PS7_RREADY;
    wire [1:0] PS7_RRESP;
    wire PS7_RVALID;
    wire [31:0] PS7_WDATA;
    wire PS7_WREADY;
    wire [3:0] PS7_WSTRB;
    wire PS7_WVALID;

    wire [31:0] M_AXI_ARADDR;
    wire M_AXI_ARREADY;
    wire  M_AXI_ARVALID;
    wire [31:0] M_AXI_AWADDR;
    wire M_AXI_AWREADY;
    wire  M_AXI_AWVALID;
    wire  M_AXI_BREADY;
    wire [1:0] M_AXI_BRESP;
    wire M_AXI_BVALID;
    wire [63:0] M_AXI_RDATA;
    wire M_AXI_RREADY;
    wire [1:0] M_AXI_RRESP;
    wire M_AXI_RVALID;
    wire [63:0] M_AXI_WDATA;
    wire M_AXI_WREADY;
    wire [7:0] M_AXI_WSTRB;
    wire M_AXI_WVALID;
    wire M_AXI_RLAST;
    wire M_AXI_WLAST;
    
    wire [3:0] M_AXI_ARLEN;
    wire [1:0] M_AXI_ARSIZE;
    wire [1:0] M_AXI_ARBURST;
    
    wire [3:0] M_AXI_AWLEN;
    wire [1:0] M_AXI_AWSIZE;
    wire [1:0] M_AXI_AWBURST;
    
    wire CONFIG_VALID;
    wire [31:0] CONFIG_CMD;
    wire [31:0] CONFIG_SRC;
    wire [31:0] CONFIG_DEST;
    wire [31:0] CONFIG_LEN;
    wire CONFIG_IRQ;
  
    wire READER_READY;
    wire WRITER_READY;
    
    assign CONFIG_READY = READER_READY && WRITER_READY;
    
    Conf conf(
    .ACLK(FCLK0),
    .ARESETN(ARESETN),
    .S_AXI_ARADDR(PS7_ARADDR), 
    .S_AXI_ARID(PS7_ARID),  
    .S_AXI_ARREADY(PS7_ARREADY), 
    .S_AXI_ARVALID(PS7_ARVALID), 
    .S_AXI_AWADDR(PS7_AWADDR), 
    .S_AXI_AWID(PS7_AWID), 
    .S_AXI_AWREADY(PS7_AWREADY), 
    .S_AXI_AWVALID(PS7_AWVALID), 
    .S_AXI_BID(PS7_BID), 
    .S_AXI_BREADY(PS7_BREADY), 
    .S_AXI_BRESP(PS7_BRESP), 
    .S_AXI_BVALID(PS7_BVALID), 
    .S_AXI_RDATA(PS7_RDATA), 
    .S_AXI_RID(PS7_RID), 
    .S_AXI_RLAST(PS7_RLAST), 
    .S_AXI_RREADY(PS7_RREADY), 
    .S_AXI_RRESP(PS7_RRESP), 
    .S_AXI_RVALID(PS7_RVALID), 
    .S_AXI_WDATA(PS7_WDATA), 
    .S_AXI_WREADY(PS7_WREADY), 
    .S_AXI_WSTRB(PS7_WSTRB), 
    .S_AXI_WVALID(PS7_WVALID),
    .CONFIG_VALID(CONFIG_VALID),
    .CONFIG_READY(CONFIG_READY),
    .CONFIG_CMD(CONFIG_CMD),
    .CONFIG_SRC(CONFIG_SRC),
    .CONFIG_DEST(CONFIG_DEST),
    .CONFIG_LEN(CONFIG_LEN),
    .CONFIG_IRQ(CONFIG_IRQ));

   // lengthInput/lengthOutput are in bytes
   wire [31:0] lengthInput;
   assign lengthInput = {4'b0000,CONFIG_LEN[27:0]};
   wire [31:0] lengthOutput;
   assign lengthOutput = (CONFIG_LEN[27:0] << 8'd8) >> CONFIG_LEN[31:28];

   reg [31:0]  clkcnt = 0;
//   assign LED = clkcnt[20:13];
   assign  LED = clkcnt[28:21];
   
  always @(posedge FCLK0) begin
//    if(ARESETN == 0)
//        LED <= 0;
//    else if(CONFIG_VALID)
//        LED <= {CONFIG_CMD[1:0],CONFIG_SRC[2:0],CONFIG_DEST[2:0]};
     clkcnt <= clkcnt+1;

  end

  wire [63:0] pipelineInput;
  wire       pipelineInputValid;
   
  wire [64:0] pipelineOutputPacked;
  wire [63:0] pipelineOutput;
  assign pipelineOutput = pipelineOutputPacked[63:0];   
  wire pipelineOutputValid;
  assign pipelineOutputValid = pipelineOutputPacked[64];
   
  wire       pipelineReady;
  wire      downstreamReady;

  
    
  harnessaxi  #(.INPUT_COUNT(76800),.OUTPUT_COUNT(153616)) pipeline(.CLK(FCLK0),.reset(CONFIG_READY),.ready(pipelineReady),.ready_downstream(downstreamReady),.process_input({pipelineInputValid,pipelineInput}),.process_output(pipelineOutputPacked));

//   UnderflowShim #(.WAIT_CYCLES(77824)) OS(.CLK(FCLK0),.RST(CONFIG_READY),.lengthOutput(lengthOutput),.inp(pipelineOutputPacked[63:0]),.inp_valid(pipelineOutputPacked[64]),.out(pipelineOutput),.out_valid(pipelineOutputValid));
   
  DRAMReader reader(
    .ACLK(FCLK0),
    .ARESETN(ARESETN),
    .M_AXI_ARADDR(M_AXI_ARADDR),
    .M_AXI_ARREADY(M_AXI_ARREADY),
    .M_AXI_ARVALID(M_AXI_ARVALID),
    .M_AXI_RDATA(M_AXI_RDATA),
    .M_AXI_RREADY(M_AXI_RREADY),
    .M_AXI_RRESP(M_AXI_RRESP),
    .M_AXI_RVALID(M_AXI_RVALID),
    .M_AXI_RLAST(M_AXI_RLAST),
    .M_AXI_ARLEN(M_AXI_ARLEN),
    .M_AXI_ARSIZE(M_AXI_ARSIZE),
    .M_AXI_ARBURST(M_AXI_ARBURST),
    
    .CONFIG_VALID(CONFIG_VALID),
    .CONFIG_READY(READER_READY),
    .CONFIG_START_ADDR(CONFIG_SRC),
    .CONFIG_NBYTES(614400),

    .DATA_READY_DOWNSTREAM(pipelineReady),
    .DATA_VALID(pipelineInputValid),
    .DATA(pipelineInput)
  );
  
  DRAMWriter writer(
    .ACLK(FCLK0),
    .ARESETN(ARESETN),
    .M_AXI_AWADDR(M_AXI_AWADDR),
    .M_AXI_AWREADY(M_AXI_AWREADY),
    .M_AXI_AWVALID(M_AXI_AWVALID),
    .M_AXI_WDATA(M_AXI_WDATA),
    .M_AXI_WREADY(M_AXI_WREADY),
    .M_AXI_WVALID(M_AXI_WVALID),
    .M_AXI_WLAST(M_AXI_WLAST),
    .M_AXI_WSTRB(M_AXI_WSTRB),
    
    .M_AXI_BRESP(M_AXI_BRESP),
    .M_AXI_BREADY(M_AXI_BREADY),
    .M_AXI_BVALID(M_AXI_BVALID),
    
    .M_AXI_AWLEN(M_AXI_AWLEN),
    .M_AXI_AWSIZE(M_AXI_AWSIZE),
    .M_AXI_AWBURST(M_AXI_AWBURST),
    
    .CONFIG_VALID(CONFIG_VALID),
    .CONFIG_READY(WRITER_READY),
    .CONFIG_START_ADDR(CONFIG_DEST),
    .CONFIG_NBYTES(1228928),

    .DATA_READY(downstreamReady),
    .DATA_VALID(pipelineOutputValid),
    .DATA(pipelineOutput)
  );

  PS7 ps7_0(
    .DMA0DATYPE(), 	// out std_logic_vector(1 downto 0);
    .DMA0DAVALID(), 	// out std_ulogic;
    .DMA0DRREADY(), 	// out std_ulogic;
    .DMA0RSTN(), 	// out std_ulogic;
    .DMA1DATYPE(), 	// out std_logic_vector(1 downto 0);
    .DMA1DAVALID(), 	// out std_ulogic;
    .DMA1DRREADY(), 	// out std_ulogic;
    .DMA1RSTN(), 	// out std_ulogic;
    .DMA2DATYPE(), 	// out std_logic_vector(1 downto 0);
    .DMA2DAVALID(), 	// out std_ulogic;
    .DMA2DRREADY(), 	// out std_ulogic;
    .DMA2RSTN(), 	// out std_ulogic;
    .DMA3DATYPE(), 	// out std_logic_vector(1 downto 0);
    .DMA3DAVALID(), 	// out std_ulogic;
    .DMA3DRREADY(), 	// out std_ulogic;
    .DMA3RSTN(), 	// out std_ulogic;
    .EMIOCAN0PHYTX(), 	// out std_ulogic;
    .EMIOCAN1PHYTX(), 	// out std_ulogic;
    .EMIOENET0GMIITXD(), 	// out std_logic_vector(7 downto 0);
    .EMIOENET0GMIITXEN(), 	// out std_ulogic;
    .EMIOENET0GMIITXER(), 	// out std_ulogic;
    .EMIOENET0MDIOMDC(), 	// out std_ulogic;
    .EMIOENET0MDIOO(), 	// out std_ulogic;
    .EMIOENET0MDIOTN(), 	// out std_ulogic;
    .EMIOENET0PTPDELAYREQRX(), 	// out std_ulogic;
    .EMIOENET0PTPDELAYREQTX(), 	// out std_ulogic;
    .EMIOENET0PTPPDELAYREQRX(), 	// out std_ulogic;
    .EMIOENET0PTPPDELAYREQTX(), 	// out std_ulogic;
    .EMIOENET0PTPPDELAYRESPRX(), 	// out std_ulogic;
    .EMIOENET0PTPPDELAYRESPTX(), 	// out std_ulogic;
    .EMIOENET0PTPSYNCFRAMERX(), 	// out std_ulogic;
    .EMIOENET0PTPSYNCFRAMETX(), 	// out std_ulogic;
    .EMIOENET0SOFRX(), 	// out std_ulogic;
    .EMIOENET0SOFTX(), 	// out std_ulogic;
    .EMIOENET1GMIITXD(), 	// out std_logic_vector(7 downto 0);
    .EMIOENET1GMIITXEN(), 	// out std_ulogic;
    .EMIOENET1GMIITXER(), 	// out std_ulogic;
    .EMIOENET1MDIOMDC(), 	// out std_ulogic;
    .EMIOENET1MDIOO(), 	// out std_ulogic;
    .EMIOENET1MDIOTN(), 	// out std_ulogic;
    .EMIOENET1PTPDELAYREQRX(), 	// out std_ulogic;
    .EMIOENET1PTPDELAYREQTX(), 	// out std_ulogic;
    .EMIOENET1PTPPDELAYREQRX(), 	// out std_ulogic;
    .EMIOENET1PTPPDELAYREQTX(), 	// out std_ulogic;
    .EMIOENET1PTPPDELAYRESPRX(), 	// out std_ulogic;
    .EMIOENET1PTPPDELAYRESPTX(), 	// out std_ulogic;
    .EMIOENET1PTPSYNCFRAMERX(), 	// out std_ulogic;
    .EMIOENET1PTPSYNCFRAMETX(), 	// out std_ulogic;
    .EMIOENET1SOFRX(), 	// out std_ulogic;
    .EMIOENET1SOFTX(), 	// out std_ulogic;
    .EMIOGPIOO(), 	 // out std_logic_vector(63 downto 0);
    .EMIOGPIOTN(),  // out std_logic_vector(63 downto 0);
    .EMIOI2C0SCLO(), 	 // out std_ulogic;
    .EMIOI2C0SCLTN(),  // out std_ulogic;
    .EMIOI2C0SDAO(), 	 // out std_ulogic;
    .EMIOI2C0SDATN(),  // out std_ulogic;
    .EMIOI2C1SCLO(), 	 // out std_ulogic;
    .EMIOI2C1SCLTN(),  // out std_ulogic;
    .EMIOI2C1SDAO(), 	 // out std_ulogic;
    .EMIOI2C1SDATN(),  // out std_ulogic;
    .EMIOPJTAGTDO(), 	// out std_ulogic;
    .EMIOPJTAGTDTN(), 	// out std_ulogic;
    .EMIOSDIO0BUSPOW(), 	// out std_ulogic;
    .EMIOSDIO0BUSVOLT(), 	// out std_logic_vector(2 downto 0);
    .EMIOSDIO0CLK(), 	// out std_ulogic;
    .EMIOSDIO0CMDO(), 	// out std_ulogic;
    .EMIOSDIO0CMDTN(), 	// out std_ulogic;
    .EMIOSDIO0DATAO(), 	// out std_logic_vector(3 downto 0);
    .EMIOSDIO0DATATN(), 	// out std_logic_vector(3 downto 0);
    .EMIOSDIO0LED(), 	// out std_ulogic;
    .EMIOSDIO1BUSPOW(), 	// out std_ulogic;
    .EMIOSDIO1BUSVOLT(), 	// out std_logic_vector(2 downto 0);
    .EMIOSDIO1CLK(), 	// out std_ulogic;
    .EMIOSDIO1CMDO(), 	// out std_ulogic;
    .EMIOSDIO1CMDTN(), 	// out std_ulogic;
    .EMIOSDIO1DATAO(), 	// out std_logic_vector(3 downto 0);
    .EMIOSDIO1DATATN(), 	// out std_logic_vector(3 downto 0);
    .EMIOSDIO1LED(), 	// out std_ulogic;
    .EMIOSPI0MO(), 	// out std_ulogic;
    .EMIOSPI0MOTN(), 	// out std_ulogic;
    .EMIOSPI0SCLKO(), 	// out std_ulogic;
    .EMIOSPI0SCLKTN(), 	// out std_ulogic;
    .EMIOSPI0SO(), 	// out std_ulogic;
    .EMIOSPI0SSNTN(), 	// out std_ulogic;
    .EMIOSPI0SSON(), 	// out std_logic_vector(2 downto 0);
    .EMIOSPI0STN(), 	// out std_ulogic;
    .EMIOSPI1MO(), 	// out std_ulogic;
    .EMIOSPI1MOTN(), 	// out std_ulogic;
    .EMIOSPI1SCLKO(), 	// out std_ulogic;
    .EMIOSPI1SCLKTN(), 	// out std_ulogic;
    .EMIOSPI1SO(), 	// out std_ulogic;
    .EMIOSPI1SSNTN(), 	// out std_ulogic;
    .EMIOSPI1SSON(), 	// out std_logic_vector(2 downto 0);
    .EMIOSPI1STN(), 	// out std_ulogic;
    .EMIOTRACECTL(), 	// out std_ulogic;
    .EMIOTRACEDATA(), 	// out std_logic_vector(31 downto 0);
    .EMIOTTC0WAVEO(), 	// out std_logic_vector(2 downto 0);
    .EMIOTTC1WAVEO(), 	// out std_logic_vector(2 downto 0);
    .EMIOUART0DTRN(), 	// out std_ulogic;
    .EMIOUART0RTSN(), 	// out std_ulogic;
    .EMIOUART0TX(), 	// out std_ulogic;
    .EMIOUART1DTRN(), 	// out std_ulogic;
    .EMIOUART1RTSN(), 	// out std_ulogic;
    .EMIOUART1TX(), 	// out std_ulogic;
    .EMIOUSB0PORTINDCTL(), 	// out std_logic_vector(1 downto 0);
    .EMIOUSB0VBUSPWRSELECT(), 	// out std_ulogic;
    .EMIOUSB1PORTINDCTL(), 	// out std_logic_vector(1 downto 0);
    .EMIOUSB1VBUSPWRSELECT(), 	// out std_ulogic;
    .EMIOWDTRSTO(), 	// out std_ulogic;
    .EVENTEVENTO(), 	// out std_ulogic;
    .EVENTSTANDBYWFE(), 	// out std_logic_vector(1 downto 0);
    .EVENTSTANDBYWFI(), 	// out std_logic_vector(1 downto 0);
    .FCLKCLK(fclk), 	 // out std_logic_vector(3 downto 0);
    .FCLKRESETN(fclkresetn), 	// out std_logic_vector(3 downto 0);
    .FTMTF2PTRIGACK(), 	// out std_logic_vector(3 downto 0);
    .FTMTP2FDEBUG(), 	// out std_logic_vector(31 downto 0);
    .FTMTP2FTRIG(), 	// out std_logic_vector(3 downto 0);
    .IRQP2F(), 	// out std_logic_vector(28 downto 0);
    
    .MAXIGP0ACLK(FCLK0), 	// in std_ulogic;
    .MAXIGP0ARADDR(PS7_ARADDR),  // out std_logic_vector(31 downto 0);
    .MAXIGP0ARBURST(),  // out std_logic_vector(1 downto 0);
    .MAXIGP0ARCACHE(),  // out std_logic_vector(3 downto 0);
    .MAXIGP0ARESETN(),  // out std_ulogic;
    .MAXIGP0ARID(PS7_ARID), 	 // out std_logic_vector(11 downto 0);
    .MAXIGP0ARLEN(),  // out std_logic_vector(3 downto 0);
    .MAXIGP0ARLOCK(),  // out std_logic_vector(1 downto 0);
    .MAXIGP0ARPROT(),  // out std_logic_vector(2 downto 0);
    .MAXIGP0ARQOS(),  // out std_logic_vector(3 downto 0);
    .MAXIGP0ARREADY(PS7_ARREADY), // in std_ulogic;
    .MAXIGP0ARSIZE(),  // out std_logic_vector(1 downto 0);
    .MAXIGP0ARVALID(PS7_ARVALID),  // out std_ulogic;
    .MAXIGP0AWADDR(PS7_AWADDR),  // out std_logic_vector(31 downto 0);
    .MAXIGP0AWBURST(),  // out std_logic_vector(1 downto 0);
    .MAXIGP0AWCACHE(),  // out std_logic_vector(3 downto 0);
    .MAXIGP0AWID(PS7_AWID), 	 // out std_logic_vector(11 downto 0);
    .MAXIGP0AWLEN(),  // out std_logic_vector(3 downto 0);
    .MAXIGP0AWLOCK(),  // out std_logic_vector(1 downto 0);
    .MAXIGP0AWPROT(),  // out std_logic_vector(2 downto 0);
    .MAXIGP0AWQOS(),  // out std_logic_vector(3 downto 0);
    .MAXIGP0AWREADY(PS7_AWREADY), // in std_ulogic;
    .MAXIGP0AWSIZE(),  // out std_logic_vector(1 downto 0);
    .MAXIGP0AWVALID(PS7_AWVALID),  // out std_ulogic;
    .MAXIGP0BID(PS7_BID), 	// in std_logic_vector(11 downto 0);
    .MAXIGP0BREADY(PS7_BREADY),  // out std_ulogic;
    .MAXIGP0BRESP(PS7_BRESP), // in std_logic_vector(1 downto 0);
    .MAXIGP0BVALID(PS7_BVALID), // in std_ulogic;
    .MAXIGP0RDATA(PS7_RDATA), // in std_logic_vector(31 downto 0);
    .MAXIGP0RID(PS7_RID), 	// in std_logic_vector(11 downto 0);
    .MAXIGP0RLAST(PS7_RLAST), // in std_ulogic;
    .MAXIGP0RREADY(PS7_RREADY),  // out std_ulogic;
    .MAXIGP0RRESP(PS7_RRESP), // in std_logic_vector(1 downto 0);    
    .MAXIGP0RVALID(PS7_RVALID), // in std_ulogic;
    .MAXIGP0WDATA(PS7_WDATA),  // out std_logic_vector(31 downto 0);
    .MAXIGP0WID(), 	 // out std_logic_vector(11 downto 0);
    .MAXIGP0WLAST(),  // out std_ulogic;
    .MAXIGP0WREADY(PS7_WREADY), // in std_ulogic;
    .MAXIGP0WSTRB(PS7_WSTRB),  // out std_logic_vector(3 downto 0);
    .MAXIGP0WVALID(PS7_WVALID),  // out std_ulogic;
    
    .MAXIGP1ARADDR(),  // out std_logic_vector(31 downto 0);
    .MAXIGP1ARBURST(),  // out std_logic_vector(1 downto 0);
    .MAXIGP1ARCACHE(),  // out std_logic_vector(3 downto 0);
    .MAXIGP1ARESETN(),  // out std_ulogic;
    .MAXIGP1ARID(), 	 // out std_logic_vector(11 downto 0);
    .MAXIGP1ARLEN(),  // out std_logic_vector(3 downto 0);
    .MAXIGP1ARLOCK(),  // out std_logic_vector(1 downto 0);
    .MAXIGP1ARPROT(),  // out std_logic_vector(2 downto 0);
    .MAXIGP1ARQOS(),  // out std_logic_vector(3 downto 0);
    .MAXIGP1ARSIZE(),  // out std_logic_vector(1 downto 0);
    .MAXIGP1ARVALID(),  // out std_ulogic;
    .MAXIGP1AWADDR(),  // out std_logic_vector(31 downto 0);
    .MAXIGP1AWBURST(),  // out std_logic_vector(1 downto 0);
    .MAXIGP1AWCACHE(),  // out std_logic_vector(3 downto 0);
    .MAXIGP1AWID(), 	 // out std_logic_vector(11 downto 0);
    .MAXIGP1AWLEN(),  // out std_logic_vector(3 downto 0);
    .MAXIGP1AWLOCK(),  // out std_logic_vector(1 downto 0);
    .MAXIGP1AWPROT(),  // out std_logic_vector(2 downto 0);
    .MAXIGP1AWQOS(),  // out std_logic_vector(3 downto 0);
    .MAXIGP1AWSIZE(),  // out std_logic_vector(1 downto 0);
    .MAXIGP1AWVALID(),  // out std_ulogic;
    .MAXIGP1BREADY(),  // out std_ulogic;
    .MAXIGP1RREADY(),  // out std_ulogic;
    .MAXIGP1WDATA(),  // out std_logic_vector(31 downto 0);
    .MAXIGP1WID(), 	 // out std_logic_vector(11 downto 0);
    .MAXIGP1WLAST(),  // out std_ulogic;
    .MAXIGP1WSTRB(),  // out std_logic_vector(3 downto 0);
    .MAXIGP1WVALID(),  // out std_ulogic;
    .SAXIGP0ARESETN(), 	// out std_ulogic;
    .SAXIGP0ARREADY(), 	// out std_ulogic;
    .SAXIGP0AWREADY(), 	// out std_ulogic;
    .SAXIGP0BID(), 	// out std_logic_vector(5 downto 0);
    .SAXIGP0BRESP(), 	// out std_logic_vector(1 downto 0);
    .SAXIGP0BVALID(), 	// out std_ulogic;
    .SAXIGP0RDATA(), 	// out std_logic_vector(31 downto 0);
    .SAXIGP0RID(), 	// out std_logic_vector(5 downto 0);
    .SAXIGP0RLAST(), 	// out std_ulogic;
    .SAXIGP0RRESP(), 	// out std_logic_vector(1 downto 0);
    .SAXIGP0RVALID(), 	// out std_ulogic;
    .SAXIGP0WREADY(), 	// out std_ulogic;
    .SAXIGP1ARESETN(), 	// out std_ulogic;
    .SAXIGP1ARREADY(), 	// out std_ulogic;
    .SAXIGP1AWREADY(), 	// out std_ulogic;
    .SAXIGP1BID(), 	// out std_logic_vector(5 downto 0);
    .SAXIGP1BRESP(), 	// out std_logic_vector(1 downto 0);
    .SAXIGP1BVALID(), 	// out std_ulogic;
    .SAXIGP1RDATA(), 	// out std_logic_vector(31 downto 0);
    .SAXIGP1RID(), 	// out std_logic_vector(5 downto 0);
    .SAXIGP1RLAST(), 	// out std_ulogic;
    .SAXIGP1RRESP(), 	// out std_logic_vector(1 downto 0);
    .SAXIGP1RVALID(), 	// out std_ulogic;
    .SAXIGP1WREADY(), 	// out std_ulogic;
    
    
    
    .SAXIHP0ACLK(1'b0), 		// in std_ulogic;
    .SAXIHP0ARADDR(32'b0),	// in std_logic_vector(31 downto 0);
    .SAXIHP0ARBURST(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIHP0ARCACHE(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIHP0ARESETN(), 	// out std_ulogic;
    .SAXIHP0ARID(6'b0),	// in std_logic_vector(2 downto 0);
    .SAXIHP0ARLEN(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIHP0ARLOCK(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIHP0ARPROT(3'b0),	// in std_logic_vector(2 downto 0);
    .SAXIHP0ARQOS(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIHP0ARREADY(), 	// out std_ulogic;
    .SAXIHP0ARSIZE(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIHP0ARVALID(1'b0), 		// in std_ulogic;
    .SAXIHP0AWADDR(32'b0),	// in std_logic_vector(31 downto 0);
    .SAXIHP0AWBURST(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIHP0AWCACHE(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIHP0AWID(6'b0),	// in std_logic_vector(2 downto 0);
    .SAXIHP0AWLEN(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIHP0AWLOCK(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIHP0AWPROT(3'b0),	// in std_logic_vector(2 downto 0);
    .SAXIHP0AWQOS(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIHP0AWREADY(), 	// out std_ulogic;
    .SAXIHP0AWSIZE(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIHP0AWVALID(1'b0), 		// in std_ulogic;
    .SAXIHP0BID(), 	// out std_logic_vector(2 downto 0);
    .SAXIHP0BREADY(1'b0), 		// in std_ulogic;
    .SAXIHP0BRESP(), 	// out std_logic_vector(1 downto 0);
    .SAXIHP0BVALID(), 	// out std_ulogic;
    .SAXIHP0RDATA(), 	// out std_logic_vector(63 downto 0);
    .SAXIHP0RID(), 	// out std_logic_vector(2 downto 0);
    .SAXIHP0RLAST(), 	// out std_ulogic;
    .SAXIHP0RREADY(1'b0), 		// in std_ulogic;
    .SAXIHP0RRESP(), 	// out std_logic_vector(1 downto 0);
    .SAXIHP0RVALID(), 	// out std_ulogic;
    .SAXIHP0WDATA(64'b0),	// in std_logic_vector(63 downto 0);
    .SAXIHP0WID(6'b0),	// in std_logic_vector(2 downto 0);
    .SAXIHP0WLAST(1'b0), 		// in std_ulogic;
    .SAXIHP0WREADY(), 	// out std_ulogic;
    .SAXIHP0WSTRB(8'b0),	// in std_logic_vector(7 downto 0);
    .SAXIHP0WVALID(1'b0), 		// in std_ulogic;
    
    .SAXIACPARUSER(5'b0),	// in std_logic_vector(4 downto 0);
    .SAXIACPAWUSER(5'b0),	// in std_logic_vector(4 downto 0);
    
    .SAXIACPACLK(FCLK0), 	// in std_ulogic;
    .SAXIACPARADDR(M_AXI_ARADDR),
    .SAXIACPARBURST(M_AXI_ARBURST), // in std_logic_vector(1 downto 0);
    .SAXIACPARCACHE(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIACPARESETN(),  // out std_ulogic;
    .SAXIACPARID(3'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIACPARLEN(M_AXI_ARLEN), // in std_logic_vector(3 downto 0);
    .SAXIACPARLOCK(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIACPARPROT(3'b0), // in std_logic_vector(2 downto 0);
    .SAXIACPARQOS(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIACPARREADY(M_AXI_ARREADY),
    .SAXIACPARSIZE(M_AXI_ARSIZE), // in std_logic_vector(1 downto 0);
    .SAXIACPARVALID(M_AXI_ARVALID),
    .SAXIACPAWADDR(M_AXI_AWADDR),
    .SAXIACPAWBURST(M_AXI_AWBURST), // in std_logic_vector(1 downto 0);
    .SAXIACPAWCACHE(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIACPAWID(3'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIACPAWLEN(M_AXI_AWLEN), // in std_logic_vector(3 downto 0);
    .SAXIACPAWLOCK(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIACPAWPROT(3'b0), // in std_logic_vector(2 downto 0);
    .SAXIACPAWQOS(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIACPAWREADY(M_AXI_AWREADY),
    .SAXIACPAWSIZE(M_AXI_AWSIZE), // in std_logic_vector(1 downto 0);
    .SAXIACPAWVALID(M_AXI_AWVALID),
    .SAXIACPBID(), 	 // out std_logic_vector(5 downto 0);
    .SAXIACPBREADY(M_AXI_BREADY),
    .SAXIACPBRESP(M_AXI_BRESP),
    .SAXIACPBVALID(M_AXI_BVALID),
    .SAXIACPRDATA(M_AXI_RDATA),
    .SAXIACPRID(), 	 // out std_logic_vector(5 downto 0);
    .SAXIACPRLAST(M_AXI_RLAST),  // out std_ulogic;
    .SAXIACPRREADY(M_AXI_RREADY),
    .SAXIACPRRESP(M_AXI_RRESP),
    .SAXIACPRVALID(M_AXI_RVALID),
    .SAXIACPWDATA(M_AXI_WDATA),
    .SAXIACPWID(3'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIACPWLAST(M_AXI_WLAST), // in std_ulogic;
    .SAXIACPWREADY(M_AXI_WREADY),
    .SAXIACPWSTRB(M_AXI_WSTRB),
    .SAXIACPWVALID(M_AXI_WVALID),
    
    .SAXIHP0RDISSUECAP1EN(1'b0), 		// in std_ulogic;
    .SAXIHP0WRISSUECAP1EN(1'b0), 		// in std_ulogic;
    .SAXIHP0RACOUNT(),  // out std_logic_vector(2 downto 0);
    .SAXIHP0RCOUNT(),  // out std_logic_vector(7 downto 0);
    .SAXIHP0WACOUNT(),  // out std_logic_vector(5 downto 0);
    .SAXIHP0WCOUNT(),  // out std_logic_vector(7 downto 0);
    
    .SAXIHP1ARESETN(),  // out std_ulogic;
    .SAXIHP1ARREADY(),  // out std_ulogic;
    .SAXIHP1AWREADY(),  // out std_ulogic;
    .SAXIHP1BID(), 	 // out std_logic_vector(5 downto 0);
    .SAXIHP1BRESP(),  // out std_logic_vector(1 downto 0);
    .SAXIHP1BVALID(),  // out std_ulogic;
    .SAXIHP1RACOUNT(),  // out std_logic_vector(2 downto 0);
    .SAXIHP1RCOUNT(),  // out std_logic_vector(7 downto 0);
    .SAXIHP1RDATA(),  // out std_logic_vector(63 downto 0);
    .SAXIHP1RID(), 	 // out std_logic_vector(5 downto 0);
    .SAXIHP1RLAST(),  // out std_ulogic;
    .SAXIHP1RRESP(),  // out std_logic_vector(1 downto 0);
    .SAXIHP1RVALID(),  // out std_ulogic;
    .SAXIHP1WACOUNT(),  // out std_logic_vector(5 downto 0);
    .SAXIHP1WCOUNT(),  // out std_logic_vector(7 downto 0);
    .SAXIHP1WREADY(),  // out std_ulogic;
    .SAXIHP2ARESETN(),  // out std_ulogic;
    .SAXIHP2ARREADY(),  // out std_ulogic;
    .SAXIHP2AWREADY(),  // out std_ulogic;
    .SAXIHP2BID(), 	 // out std_logic_vector(5 downto 0);
    .SAXIHP2BRESP(),  // out std_logic_vector(1 downto 0);
    .SAXIHP2BVALID(),  // out std_ulogic;
    .SAXIHP2RACOUNT(),  // out std_logic_vector(2 downto 0);
    .SAXIHP2RCOUNT(),  // out std_logic_vector(7 downto 0);
    .SAXIHP2RDATA(),  // out std_logic_vector(63 downto 0);
    .SAXIHP2RID(), 	 // out std_logic_vector(5 downto 0);
    .SAXIHP2RLAST(),  // out std_ulogic;
    .SAXIHP2RRESP(),  // out std_logic_vector(1 downto 0);
    .SAXIHP2RVALID(),  // out std_ulogic;
    .SAXIHP2WACOUNT(),  // out std_logic_vector(5 downto 0);
    .SAXIHP2WCOUNT(),  // out std_logic_vector(7 downto 0);
    .SAXIHP2WREADY(),  // out std_ulogic;
    .SAXIHP3ARESETN(),  // out std_ulogic;
    .SAXIHP3ARREADY(),  // out std_ulogic;
    .SAXIHP3AWREADY(),  // out std_ulogic;
    .SAXIHP3BID(), 	 // out std_logic_vector(5 downto 0);
    .SAXIHP3BRESP(),  // out std_logic_vector(1 downto 0);
    .SAXIHP3BVALID(),  // out std_ulogic;
    .SAXIHP3RACOUNT(),  // out std_logic_vector(2 downto 0);
    .SAXIHP3RCOUNT(),  // out std_logic_vector(7 downto 0);
    .SAXIHP3RDATA(),  // out std_logic_vector(63 downto 0);
    .SAXIHP3RID(), 	 // out std_logic_vector(5 downto 0);
    .SAXIHP3RLAST(),  // out std_ulogic;
    .SAXIHP3RRESP(),  // out std_logic_vector(1 downto 0);
    .SAXIHP3RVALID(),  // out std_ulogic;
    .SAXIHP3WACOUNT(),  // out std_logic_vector(5 downto 0);
    .SAXIHP3WCOUNT(),  // out std_logic_vector(7 downto 0);
    .SAXIHP3WREADY(),  // out std_ulogic;
    .DDRA(DDR_Addr), 	// inout std_logic_vector(14 downto 0);
    .DDRBA(DDR_BankAddr), // inout std_logic_vector(2 downto 0);
    .DDRCASB(DDR_CAS_n), 	// inout std_ulogic;
    .DDRCKE(DDR_CKE), 	// inout std_ulogic;
    .DDRCKN(DDR_Clk_n), 	// inout std_ulogic;
    .DDRCKP(DDR_Clk), 	// inout std_ulogic;
    .DDRCSB(DDR_CS_n), 	// inout std_ulogic;
    .DDRDM(DDR_DM), 	// inout std_logic_vector(3 downto 0);
    .DDRDQ(DDR_DQ), 	// inout std_logic_vector(31 downto 0);
    .DDRDQSN(DDR_DQS_n), 	// inout std_logic_vector(3 downto 0);
    .DDRDQSP(DDR_DQS), 	// inout std_logic_vector(3 downto 0);
    .DDRDRSTB(DDR_DRSTB), 	// inout std_ulogic;
    .DDRODT(DDR_ODT), 	// inout std_ulogic;
    .DDRRASB(DDR_RAS_n), 	// inout std_ulogic;
    .DDRVRN(DDR_VRN), 	// inout std_ulogic;
    .DDRVRP(DDR_VRP), 	// inout std_ulogic;
    .DDRWEB(DDR_WEB), 	// inout std_ulogic;
    .MIO(MIO), 	// inout std_logic_vector(53 downto 0);
    .PSCLK(PS_CLK), 	// inout std_ulogic;
    .PSPORB(PS_PORB), 	// inout std_ulogic;
    .PSSRSTB(PS_SRSTB), 	// inout std_ulogic;
    .DDRARB(4'b0),	// in std_logic_vector(3 downto 0);
    .DMA0ACLK(1'b0), 		// in std_ulogic;
    .DMA0DAREADY(1'b0), 		// in std_ulogic;
    .DMA0DRLAST(1'b0), 		// in std_ulogic;
    .DMA0DRTYPE(2'b0),	// in std_logic_vector(1 downto 0);
    .DMA0DRVALID(1'b0), 		// in std_ulogic;
    .DMA1ACLK(1'b0), 		// in std_ulogic;
    .DMA1DAREADY(1'b0), 		// in std_ulogic;
    .DMA1DRLAST(1'b0), 		// in std_ulogic;
    .DMA1DRTYPE(2'b0),	// in std_logic_vector(1 downto 0);
    .DMA1DRVALID(1'b0), 		// in std_ulogic;
    .DMA2ACLK(1'b0), 		// in std_ulogic;
    .DMA2DAREADY(1'b0), 		// in std_ulogic;
    .DMA2DRLAST(1'b0), 		// in std_ulogic;
    .DMA2DRTYPE(2'b0),	// in std_logic_vector(1 downto 0);
    .DMA2DRVALID(1'b0), 		// in std_ulogic;
    .DMA3ACLK(1'b0), 		// in std_ulogic;
    .DMA3DAREADY(1'b0), 		// in std_ulogic;
    .DMA3DRLAST(1'b0), 		// in std_ulogic;
    .DMA3DRTYPE(2'b0),	// in std_logic_vector(1 downto 0);
    .DMA3DRVALID(1'b0), 		// in std_ulogic;
    .EMIOCAN0PHYRX(1'b0), 		// in std_ulogic;
    .EMIOCAN1PHYRX(1'b0), 		// in std_ulogic;
    .EMIOENET0EXTINTIN(1'b0), 		// in std_ulogic;
    .EMIOENET0GMIICOL(1'b0), 		// in std_ulogic;
    .EMIOENET0GMIICRS(1'b0), 		// in std_ulogic;
    .EMIOENET0GMIIRXCLK(1'b0), 		// in std_ulogic;
    .EMIOENET0GMIIRXD(8'b0),	// in std_logic_vector(7 downto 0);
    .EMIOENET0GMIIRXDV(1'b0), 		// in std_ulogic;
    .EMIOENET0GMIIRXER(1'b0), 		// in std_ulogic;
    .EMIOENET0GMIITXCLK(1'b0), 		// in std_ulogic;
    .EMIOENET0MDIOI(1'b0), 		// in std_ulogic;
    .EMIOENET1EXTINTIN(1'b0), 		// in std_ulogic;
    .EMIOENET1GMIICOL(1'b0), 		// in std_ulogic;
    .EMIOENET1GMIICRS(1'b0), 		// in std_ulogic;
    .EMIOENET1GMIIRXCLK(1'b0), 		// in std_ulogic;
    .EMIOENET1GMIIRXD(8'b0),	// in std_logic_vector(7 downto 0);
    .EMIOENET1GMIIRXDV(1'b0), 		// in std_ulogic;
    .EMIOENET1GMIIRXER(1'b0), 		// in std_ulogic;
    .EMIOENET1GMIITXCLK(1'b0), 		// in std_ulogic;
    .EMIOENET1MDIOI(1'b0), 		// in std_ulogic;
    .EMIOGPIOI(64'b0), 	// in std_logic_vector(63 downto 0);
    .EMIOI2C0SCLI(1'b0), 	// in std_ulogic;
    .EMIOI2C0SDAI(1'b0), 	// in std_ulogic;
    .EMIOI2C1SCLI(1'b0), 	// in std_ulogic;
    .EMIOI2C1SDAI(1'b0), 	// in std_ulogic;
    .EMIOPJTAGTCK(1'b0), 		// in std_ulogic;
    .EMIOPJTAGTDI(1'b0), 		// in std_ulogic;
    .EMIOPJTAGTMS(1'b0), 		// in std_ulogic;
    .EMIOSDIO0CDN(1'b0), 		// in std_ulogic;
    .EMIOSDIO0CLKFB(1'b0), 		// in std_ulogic;
    .EMIOSDIO0CMDI(1'b0), 		// in std_ulogic;
    .EMIOSDIO0DATAI(4'b0),	// in std_logic_vector(3 downto 0);
    .EMIOSDIO0WP(1'b0), 		// in std_ulogic;
    .EMIOSDIO1CDN(1'b0), 		// in std_ulogic;
    .EMIOSDIO1CLKFB(1'b0), 		// in std_ulogic;
    .EMIOSDIO1CMDI(1'b0), 		// in std_ulogic;
    .EMIOSDIO1DATAI(4'b0),	// in std_logic_vector(3 downto 0);
    .EMIOSDIO1WP(1'b0), 		// in std_ulogic;
    .EMIOSPI0MI(1'b0), 		// in std_ulogic;
    .EMIOSPI0SCLKI(1'b0), 		// in std_ulogic;
    .EMIOSPI0SI(1'b0), 		// in std_ulogic;
    .EMIOSPI0SSIN(1'b0), 		// in std_ulogic;
    .EMIOSPI1MI(1'b0), 		// in std_ulogic;
    .EMIOSPI1SCLKI(1'b0), 		// in std_ulogic;
    .EMIOSPI1SI(1'b0), 		// in std_ulogic;
    .EMIOSPI1SSIN(1'b0), 		// in std_ulogic;
    .EMIOSRAMINTIN(1'b0), 		// in std_ulogic;
    .EMIOTRACECLK(1'b0), 		// in std_ulogic;
    .EMIOTTC0CLKI(3'b0),	// in std_logic_vector(2 downto 0);
    .EMIOTTC1CLKI(3'b0),	// in std_logic_vector(2 downto 0);
    .EMIOUART0CTSN(1'b0), 		// in std_ulogic;
    .EMIOUART0DCDN(1'b0), 		// in std_ulogic;
    .EMIOUART0DSRN(1'b0), 		// in std_ulogic;
    .EMIOUART0RIN(1'b0), 		// in std_ulogic;
    .EMIOUART0RX(1'b0), 		// in std_ulogic;
    .EMIOUART1CTSN(1'b0), 		// in std_ulogic;
    .EMIOUART1DCDN(1'b0), 		// in std_ulogic;
    .EMIOUART1DSRN(1'b0), 		// in std_ulogic;
    .EMIOUART1RIN(1'b0), 		// in std_ulogic;
    .EMIOUART1RX(1'b0), 		// in std_ulogic;
    .EMIOUSB0VBUSPWRFAULT(1'b0), 		// in std_ulogic;
    .EMIOUSB1VBUSPWRFAULT(1'b0), 		// in std_ulogic;
    .EMIOWDTCLKI(1'b0), 		// in std_ulogic;
    .EVENTEVENTI(1'b0), 		// in std_ulogic;
    .FCLKCLKTRIGN(4'b0),	// in std_logic_vector(3 downto 0);
    .FPGAIDLEN(1'b0), 		// in std_ulogic;
    .FTMDTRACEINATID(4'b0),	// in std_logic_vector(3 downto 0);
    .FTMDTRACEINCLOCK(1'b0), 		// in std_ulogic;
    .FTMDTRACEINDATA(32'b0),	// in std_logic_vector(31 downto 0);
    .FTMDTRACEINVALID(1'b0), 		// in std_ulogic;
    .FTMTF2PDEBUG(32'b0),	// in std_logic_vector(31 downto 0);
    .FTMTF2PTRIG(4'b0),	// in std_logic_vector(3 downto 0);
    .FTMTP2FTRIGACK(4'b0),	// in std_logic_vector(3 downto 0);
    .IRQF2P({19'b0,CONFIG_IRQ}),	// in std_logic_vector(19 downto 0);
    .MAXIGP1ACLK(1'b0), 	// in std_ulogic;
    .MAXIGP1ARREADY(1'b0), // in std_ulogic;
    .MAXIGP1AWREADY(1'b0), // in std_ulogic;
    .MAXIGP1BID(12'b0), 	// in std_logic_vector(11 downto 0);
    .MAXIGP1BRESP(2'b0), // in std_logic_vector(1 downto 0);
    .MAXIGP1BVALID(1'b0), // in std_ulogic;
    .MAXIGP1RDATA(32'b0), // in std_logic_vector(31 downto 0);
    .MAXIGP1RID(12'b0), 	// in std_logic_vector(11 downto 0);
    .MAXIGP1RLAST(1'b0), // in std_ulogic;
    .MAXIGP1RRESP(2'b0), // in std_logic_vector(1 downto 0);
    .MAXIGP1RVALID(1'b0), // in std_ulogic;
    .MAXIGP1WREADY(1'b0), // in std_ulogic;
    .SAXIGP0ACLK(1'b0), 		// in std_ulogic;
    .SAXIGP0ARADDR(32'b0),	// in std_logic_vector(31 downto 0);
    .SAXIGP0ARBURST(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP0ARCACHE(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP0ARID(6'b0),	// in std_logic_vector(5 downto 0);
    .SAXIGP0ARLEN(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP0ARLOCK(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP0ARPROT(3'b0),	// in std_logic_vector(2 downto 0);
    .SAXIGP0ARQOS(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP0ARSIZE(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP0ARVALID(1'b0), 		// in std_ulogic;
    .SAXIGP0AWADDR(32'b0),	// in std_logic_vector(31 downto 0);
    .SAXIGP0AWBURST(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP0AWCACHE(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP0AWID(6'b0),	// in std_logic_vector(5 downto 0);
    .SAXIGP0AWLEN(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP0AWLOCK(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP0AWPROT(3'b0),	// in std_logic_vector(2 downto 0);
    .SAXIGP0AWQOS(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP0AWSIZE(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP0AWVALID(1'b0), 		// in std_ulogic;
    .SAXIGP0BREADY(1'b0), 		// in std_ulogic;
    .SAXIGP0RREADY(1'b0), 		// in std_ulogic;
    .SAXIGP0WDATA(32'b0),	// in std_logic_vector(31 downto 0);
    .SAXIGP0WID(6'b0),	// in std_logic_vector(5 downto 0);
    .SAXIGP0WLAST(1'b0), 		// in std_ulogic;
    .SAXIGP0WSTRB(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP0WVALID(1'b0), 		// in std_ulogic;
    .SAXIGP1ACLK(1'b0), 		// in std_ulogic;
    .SAXIGP1ARADDR(32'b0),	// in std_logic_vector(31 downto 0);
    .SAXIGP1ARBURST(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP1ARCACHE(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP1ARID(6'b0),	// in std_logic_vector(5 downto 0);
    .SAXIGP1ARLEN(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP1ARLOCK(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP1ARPROT(3'b0),	// in std_logic_vector(2 downto 0);
    .SAXIGP1ARQOS(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP1ARSIZE(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP1ARVALID(1'b0), 		// in std_ulogic;
    .SAXIGP1AWADDR(32'b0),	// in std_logic_vector(31 downto 0);
    .SAXIGP1AWBURST(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP1AWCACHE(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP1AWID(6'b0),	// in std_logic_vector(5 downto 0);
    .SAXIGP1AWLEN(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP1AWLOCK(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP1AWPROT(3'b0),	// in std_logic_vector(2 downto 0);
    .SAXIGP1AWQOS(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP1AWSIZE(2'b0),	// in std_logic_vector(1 downto 0);
    .SAXIGP1AWVALID(1'b0), 		// in std_ulogic;
    .SAXIGP1BREADY(1'b0), 		// in std_ulogic;
    .SAXIGP1RREADY(1'b0), 		// in std_ulogic;
    .SAXIGP1WDATA(32'b0),	// in std_logic_vector(31 downto 0);
    .SAXIGP1WID(6'b0),	// in std_logic_vector(5 downto 0);
    .SAXIGP1WLAST(1'b0), 		// in std_ulogic;
    .SAXIGP1WSTRB(4'b0),	// in std_logic_vector(3 downto 0);
    .SAXIGP1WVALID(1'b0), 		// in std_ulogic;
    .SAXIHP1ACLK(1'b0), 	// in std_ulogic;
    .SAXIHP1ARADDR(32'b0), // in std_logic_vector(31 downto 0);
    .SAXIHP1ARBURST(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP1ARCACHE(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP1ARID(6'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIHP1ARLEN(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP1ARLOCK(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP1ARPROT(3'b0), // in std_logic_vector(2 downto 0);
    .SAXIHP1ARQOS(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP1ARSIZE(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP1ARVALID(1'b0), // in std_ulogic;
    .SAXIHP1AWADDR(32'b0), // in std_logic_vector(31 downto 0);
    .SAXIHP1AWBURST(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP1AWCACHE(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP1AWID(6'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIHP1AWLEN(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP1AWLOCK(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP1AWPROT(3'b0), // in std_logic_vector(2 downto 0);
    .SAXIHP1AWQOS(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP1AWSIZE(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP1AWVALID(1'b0), // in std_ulogic;
    .SAXIHP1BREADY(1'b0), // in std_ulogic;
    .SAXIHP1RDISSUECAP1EN(1'b0), 		// in std_ulogic;
    .SAXIHP1RREADY(1'b0), // in std_ulogic;
    .SAXIHP1WDATA(64'b0), // in std_logic_vector(63 downto 0);
    .SAXIHP1WID(6'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIHP1WLAST(1'b0), // in std_ulogic;
    .SAXIHP1WRISSUECAP1EN(1'b0), 		// in std_ulogic;
    .SAXIHP1WSTRB(8'b0), // in std_logic_vector(7 downto 0);
    .SAXIHP1WVALID(1'b0), // in std_ulogic;
    .SAXIHP2ACLK(1'b0), 	// in std_ulogic;
    .SAXIHP2ARADDR(32'b0), // in std_logic_vector(31 downto 0);
    .SAXIHP2ARBURST(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP2ARCACHE(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP2ARID(6'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIHP2ARLEN(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP2ARLOCK(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP2ARPROT(3'b0), // in std_logic_vector(2 downto 0);
    .SAXIHP2ARQOS(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP2ARSIZE(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP2ARVALID(1'b0), // in std_ulogic;
    .SAXIHP2AWADDR(32'b0), // in std_logic_vector(31 downto 0);
    .SAXIHP2AWBURST(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP2AWCACHE(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP2AWID(6'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIHP2AWLEN(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP2AWLOCK(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP2AWPROT(3'b0), // in std_logic_vector(2 downto 0);
    .SAXIHP2AWQOS(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP2AWSIZE(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP2AWVALID(1'b0), // in std_ulogic;
    .SAXIHP2BREADY(1'b0), // in std_ulogic;
    .SAXIHP2RDISSUECAP1EN(1'b0), 		// in std_ulogic;
    .SAXIHP2RREADY(1'b0), // in std_ulogic;
    .SAXIHP2WDATA(64'b0), // in std_logic_vector(63 downto 0);
    .SAXIHP2WID(6'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIHP2WLAST(1'b0), // in std_ulogic;
    .SAXIHP2WRISSUECAP1EN(1'b0), 		// in std_ulogic;
    .SAXIHP2WSTRB(8'b0), // in std_logic_vector(7 downto 0);
    .SAXIHP2WVALID(1'b0), // in std_ulogic;
    .SAXIHP3ACLK(1'b0), 	// in std_ulogic;
    .SAXIHP3ARADDR(32'b0), // in std_logic_vector(31 downto 0);
    .SAXIHP3ARBURST(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP3ARCACHE(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP3ARID(6'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIHP3ARLEN(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP3ARLOCK(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP3ARPROT(3'b0), // in std_logic_vector(2 downto 0);
    .SAXIHP3ARQOS(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP3ARSIZE(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP3ARVALID(1'b0), // in std_ulogic;
    .SAXIHP3AWADDR(32'b0), // in std_logic_vector(31 downto 0);
    .SAXIHP3AWBURST(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP3AWCACHE(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP3AWID(6'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIHP3AWLEN(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP3AWLOCK(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP3AWPROT(3'b0), // in std_logic_vector(2 downto 0);
    .SAXIHP3AWQOS(4'b0), // in std_logic_vector(3 downto 0);
    .SAXIHP3AWSIZE(2'b0), // in std_logic_vector(1 downto 0);
    .SAXIHP3AWVALID(1'b0), // in std_ulogic;
    .SAXIHP3BREADY(1'b0), // in std_ulogic;
    .SAXIHP3RDISSUECAP1EN(1'b0), 		// in std_ulogic;
    .SAXIHP3RREADY(1'b0), // in std_ulogic;
    .SAXIHP3WDATA(64'b0), // in std_logic_vector(63 downto 0);
    .SAXIHP3WID(6'b0), 	// in std_logic_vector(5 downto 0);
    .SAXIHP3WLAST(1'b0), // in std_ulogic;
    .SAXIHP3WRISSUECAP1EN(1'b0), 		// in std_ulogic;
    .SAXIHP3WSTRB(8'b0), // in std_logic_vector(7 downto 0);
    .SAXIHP3WVALID(1'b0)	// in std_ulogic;
  );
endmodule
