module display(


    vga vga_inst(
        .clk_25_175_kHz(clk_25_175kHz),
        .rst_n(rst_n),
        .HS_n,
        .VS_n,
        .pixel_valid,
        .vga_row,
        .vga_col
    );


);






endmodule : display
